module dct(input [2:0] x, y, u, v, output reg [31:0] coef);
reg new_n0_, new_n1_, new_n2_, new_n3_, new_n4_, new_n5_, new_n6_, new_n7_, new_n8_, new_n9_, new_n10_, new_n11_, new_n12_, new_n13_, new_n14_, new_n15_, new_n16_, new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_;
always @(*) begin
casez ({new_n96_, new_n5848_, new_n342_, new_n3279_, new_n929_, new_n4331_, v[0], new_n5950_, new_n1257_, new_n5420_, new_n107_, new_n709_, new_n694_, new_n5111_, new_n1259_, new_n2990_, new_n109_, new_n550_, new_n883_, new_n5070_, new_n236_, new_n1090_, new_n436_, new_n6025_, new_n612_, new_n722_, new_n240_, new_n2954_, new_n121_, new_n1913_, new_n194_, new_n221_, new_n730_, new_n148_, new_n166_, new_n445_, new_n6136_, new_n1762_, new_n234_, new_n5221_, new_n122_, new_n2953_, new_n140_, new_n1370_, new_n82_, new_n154_, new_n766_})
47'b10????????????????????????????????????????????? : coef[0] = 1'b1;
47'b??11??????????????????????????????????????????? : coef[0] = 1'b1;
47'b????11????????????????????????????????????????? : coef[0] = 1'b1;
47'b??????10??????????????????????????????????????? : coef[0] = 1'b1;
47'b????????10????????????????????????????????????? : coef[0] = 1'b1;
47'b??????????00??????????????????????????????????? : coef[0] = 1'b1;
47'b????????????00????????????????????????????????? : coef[0] = 1'b1;
47'b??????????????10??????????????????????????????? : coef[0] = 1'b1;
47'b????????????????00????????????????????????????? : coef[0] = 1'b1;
47'b??????????????????01??????????????????????????? : coef[0] = 1'b1;
47'b????????????????????11????????????????????????? : coef[0] = 1'b1;
47'b??????????????????????10??????????????????????? : coef[0] = 1'b1;
47'b????????????????????????1?????????????????????? : coef[0] = 1'b1;
47'b?????????????????????????1????????????????????? : coef[0] = 1'b1;
47'b??????????????????????????11??????????????????? : coef[0] = 1'b1;
47'b????????????????????????????11????????????????? : coef[0] = 1'b1;
47'b??????????????????????????????111?????????????? : coef[0] = 1'b1;
47'b?????????????????????????????????111??????????? : coef[0] = 1'b1;
47'b??????0?????????????????????????????0?????????? : coef[0] = 1'b1;
47'b?????????????????????????????????????0????????? : coef[0] = 1'b1;
47'b??????????????????????????????????????10??????? : coef[0] = 1'b1;
47'b????????????????????????????????????????11????? : coef[0] = 1'b1;
47'b??????????????????????????????????????????11??? : coef[0] = 1'b1;
47'b????????????????????????????????????????????111 : coef[0] = 1'b1;
default : coef[0] = 1'b0;
endcase
casez ({new_n480_, new_n994_, new_n360_, new_n4687_, new_n228_, new_n419_, new_n138_, new_n5032_, new_n94_, new_n5810_, new_n339_, new_n1175_, y[1], new_n3992_, new_n2040_, new_n460_, new_n3672_, new_n398_, new_n4985_, new_n505_, new_n1180_, new_n230_, new_n1876_, new_n391_, new_n3447_, new_n2870_, new_n2567_, new_n530_, new_n1462_, new_n306_, new_n5892_, new_n716_, new_n1174_, new_n310_, new_n1652_, new_n292_, new_n3123_, new_n261_, new_n4745_, new_n667_, new_n1552_, new_n226_, new_n3329_, new_n150_, new_n2561_, new_n129_, new_n5374_, new_n101_, new_n5929_, u[0], new_n5957_, new_n1099_, new_n2770_, new_n88_, new_n696_, new_n115_, new_n3251_, new_n139_, new_n1496_, new_n425_, new_n2957_, new_n185_, new_n1019_, new_n277_, new_n1931_, new_n253_, new_n497_, new_n911_, new_n3224_, new_n301_, new_n5891_, new_n545_, new_n3282_, u[1], new_n727_, new_n222_, new_n6131_, new_n679_, new_n1765_, new_n623_, new_n3005_, new_n259_, new_n3125_, new_n818_, new_n2497_, new_n1258_, new_n3880_, new_n355_, new_n3079_, new_n224_, new_n3636_, u[2], new_n254_, new_n2851_, new_n324_, new_n5330_, new_n127_, new_n1136_, new_n299_, new_n5246_, new_n2652_, new_n5245_, new_n136_, new_n2752_, new_n183_, new_n1104_, new_n363_, new_n986_, new_n287_, new_n723_, new_n81_, new_n1832_, new_n495_, new_n1340_, new_n783_, new_n1953_, v[2], new_n3780_, new_n395_, new_n3608_, new_n493_, new_n4788_, new_n796_, new_n980_, new_n204_, new_n942_, new_n77_, new_n4798_, new_n2246_, new_n274_, new_n1473_, new_n390_, new_n578_, new_n601_, new_n712_, new_n121_, new_n948_, new_n212_, new_n649_, new_n153_, new_n908_, new_n794_, new_n1799_, new_n281_, new_n902_, new_n110_, new_n3459_, new_n113_, new_n692_, new_n172_, new_n5773_, new_n171_, new_n5485_, new_n374_, new_n3262_, new_n103_, new_n1037_, new_n80_, new_n160_, new_n2783_, new_n503_, new_n695_, new_n251_, new_n3188_, new_n137_, new_n4093_, new_n266_, new_n4877_, new_n169_, new_n1463_, new_n179_, new_n4830_, new_n404_, new_n5720_, new_n170_, new_n5588_, new_n96_, new_n5940_, new_n168_, new_n5993_, new_n269_, new_n3363_, new_n199_, new_n5211_, new_n189_, new_n4566_, new_n603_, new_n4383_, new_n557_, new_n964_, new_n300_, new_n5170_, new_n240_, new_n5949_, new_n213_, new_n1722_, new_n211_, new_n5942_, new_n284_, new_n1070_, new_n272_, new_n682_, new_n175_, new_n5719_, new_n795_, new_n4677_, new_n246_, new_n4161_, new_n196_, new_n6093_, new_n1891_, new_n4866_, new_n166_, new_n5754_, new_n219_, new_n1761_, new_n361_, new_n2759_, new_n318_, new_n5506_, new_n457_, new_n2695_, new_n167_, new_n1776_, new_n86_, new_n814_, new_n202_, new_n3708_, new_n123_, new_n5527_, new_n461_, new_n792_, new_n1902_, new_n1954_, new_n558_, new_n4648_, new_n84_, new_n87_, new_n2114_, new_n205_, new_n1178_, new_n128_, new_n4434_, new_n191_, new_n5663_, new_n248_, new_n972_, new_n354_, new_n1962_, new_n1474_, new_n2912_, new_n537_, new_n1160_, new_n868_, new_n1035_, new_n389_, new_n1385_, new_n634_, new_n4222_, new_n430_, new_n5748_, new_n273_, new_n1730_, new_n1064_, new_n2932_, new_n329_, new_n604_, new_n1620_, new_n4867_, new_n267_, new_n1585_, new_n741_, new_n3348_, new_n369_, new_n1746_, new_n1976_, new_n5439_, new_n469_, new_n5083_, new_n377_, new_n3544_, new_n2501_, new_n3799_, new_n122_, new_n5791_, new_n148_, new_n3243_, new_n371_, new_n2789_, new_n517_, new_n1228_, new_n429_, new_n1798_, new_n953_, new_n3335_, new_n455_, new_n632_, new_n262_, new_n1435_, new_n864_, new_n958_, new_n372_, new_n3721_, new_n159_, new_n860_, new_n192_, new_n643_, new_n334_, new_n5780_, new_n201_, new_n1787_, new_n1371_, new_n3092_, new_n554_, new_n1503_, new_n176_, new_n3971_, new_n869_, new_n4101_, new_n386_, new_n5961_, new_n819_, new_n1816_, new_n509_, new_n5068_, new_n733_, new_n2941_, new_n427_, new_n1617_, new_n368_, new_n5080_, new_n231_, new_n2837_, new_n642_, new_n3216_, new_n2365_, new_n311_, new_n582_, new_n375_, new_n5057_, new_n164_, new_n5969_, new_n278_, new_n4607_, new_n5432_, new_n200_, new_n1378_, new_n1171_, new_n3410_, new_n263_, new_n5963_, new_n303_, new_n1163_, new_n385_, new_n6097_, new_n151_, new_n780_, new_n332_, new_n2991_, new_n182_, new_n4345_, new_n791_, new_n1949_, new_n214_, new_n2657_, new_n223_, new_n5267_, new_n178_, new_n2819_, new_n2156_, new_n3772_, new_n85_, new_n89_, new_n782_, new_n409_, new_n751_, new_n268_, new_n1733_, new_n190_, new_n1498_, x[1], new_n187_, new_n2757_, new_n875_, new_n3591_, new_n145_, new_n745_, new_n2880_, new_n910_, new_n3141_, new_n174_, new_n5342_, new_n229_, new_n280_, new_n238_, new_n621_, new_n239_, new_n3555_})
398'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????0???????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????010???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????010?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101???????????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??????????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[1] = 1'b0;
398'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[1] = 1'b0;
398'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[1] = 1'b0;
398'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[1] = 1'b0;
398'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[1] = 1'b0;
default : coef[1] = 1'b1;
endcase
casez ({new_n648_, new_n793_, new_n360_, new_n2585_, new_n504_, new_n1752_, new_n460_, new_n1910_, new_n271_, new_n383_, new_n225_, new_n2277_, new_n442_, new_n3491_, new_n174_, new_n2673_, new_n6238_, new_n122_, new_n645_, new_n522_, new_n1050_, new_n262_, new_n4683_, new_n486_, new_n5144_, new_n2324_, new_n783_, new_n865_, new_n247_, new_n2590_, new_n121_, new_n5907_, new_n6195_, new_n1034_, new_n4418_, new_n744_, new_n1649_, new_n309_, new_n881_, new_n505_, new_n4175_, new_n633_, new_n4471_, new_n388_, new_n2829_, new_n604_, new_n678_, new_n1802_, new_n4413_, new_n191_, new_n5391_, new_n864_, new_n3600_, new_n215_, new_n5475_, new_n154_, new_n4142_, new_n317_, new_n949_, new_n447_, new_n2769_, new_n339_, new_n1848_, new_n1892_, new_n4208_, new_n86_, new_n493_, new_n1035_, new_n103_, new_n3928_, new_n251_, new_n4454_, new_n356_, new_n5263_, new_n211_, new_n2004_, new_n142_, new_n5639_, new_n153_, new_n5935_, new_n115_, new_n2723_, new_n389_, new_n669_, new_n1201_, new_n4461_, new_n2483_, new_n294_, new_n4013_, new_n1549_, new_n4145_, new_n237_, new_n4832_, new_n137_, new_n4949_, new_n168_, new_n5513_, new_n2275_, new_n131_, new_n3354_, new_n249_, new_n1059_, new_n1577_, new_n3968_, new_n285_, new_n1346_, new_n279_, new_n2797_, new_n171_, new_n5974_, new_n307_, new_n1482_, new_n2860_, new_n2859_, new_n151_, new_n843_, new_n179_, new_n5241_, new_n166_, new_n374_, new_n6228_, new_n2455_, new_n226_, new_n1694_, new_n426_, new_n2163_, new_n268_, new_n4237_, new_n521_, new_n1550_, new_n113_, new_n6192_, new_n266_, new_n758_, new_n172_, new_n762_, new_n300_, new_n6109_, new_n164_, new_n1155_, new_n269_, new_n4466_, new_n254_, new_n5496_, new_n293_, new_n3948_, new_n2809_, new_n4690_, new_n3442_, new_n313_, new_n2121_, new_n427_, new_n1490_, new_n554_, new_n4966_, new_n344_, new_n2845_, new_n746_, new_n3671_, new_n253_, new_n4203_, new_n312_, new_n5329_, new_n325_, new_n496_, new_n272_, new_n4449_, new_n186_, new_n3151_, new_n175_, new_n5520_, new_n183_, new_n1598_, new_n422_, new_n3150_, new_n157_, new_n6084_, new_n182_, new_n3774_, new_n347_, new_n612_, new_n305_, new_n2597_, new_n509_, new_n2666_, new_n982_, new_n1570_, new_n525_, new_n4349_, new_n91_, new_n1604_, new_n286_, new_n534_, new_n94_, new_n160_, new_n750_, new_n177_, new_n464_, new_n145_, new_n4509_, new_n202_, new_n635_, new_n128_, new_n3713_, new_n178_, new_n1874_, new_n241_, new_n1559_, new_n502_, new_n967_, new_n542_, new_n2770_, new_n184_, new_n1459_, new_n420_, new_n3505_, new_n161_, new_n910_, new_n155_, new_n3938_, new_n213_, new_n2615_, new_n457_, new_n4404_, new_n189_, new_n756_, new_n248_, new_n1077_, new_n5432_, new_n346_, new_n1477_, new_n673_, new_n3583_, new_n144_, new_n2094_, new_n167_, new_n880_, new_n602_, new_n1041_, new_n208_, new_n6164_, new_n1071_, new_n4551_, new_n503_, new_n697_, new_n672_, new_n3090_, new_n258_, new_n5929_, new_n500_, new_n1745_, u[1], new_n1899_, new_n263_, new_n5089_, new_n6240_, new_n129_, new_n4217_, new_n715_, new_n1543_, new_n281_, new_n1070_, new_n176_, new_n4801_, new_n950_, new_n1386_, new_n222_, new_n4382_, new_n452_, new_n5792_, new_n410_, new_n3586_, new_n159_, new_n1748_, new_n273_, new_n1475_, new_n434_, new_n2774_, new_n433_, new_n896_, new_n277_, new_n2047_, new_n239_, new_n5698_, new_n6225_, new_n229_, new_n1759_, new_n2748_, new_n3835_, new_n398_, new_n1714_, new_n582_, new_n972_, new_n812_, new_n1566_, new_n201_, new_n4741_, new_n205_, new_n1879_, new_n676_, new_n1486_, new_n199_, new_n5345_, new_n6250_})
304'b11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????? : coef[2] = 1'b1;
304'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[2] = 1'b1;
304'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??? : coef[2] = 1'b1;
304'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11? : coef[2] = 1'b1;
304'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0 : coef[2] = 1'b1;
default : coef[2] = 1'b0;
endcase
casez ({new_n487_, new_n1921_, new_n2211_, new_n486_, new_n1481_, new_n89_, new_n221_, new_n435_, new_n740_, new_n3073_, new_n176_, new_n5696_, new_n1737_, new_n2511_, new_n225_, new_n6002_, y[0], new_n1006_, new_n504_, new_n5700_, new_n283_, new_n416_, v[2], new_n215_, new_n309_, new_n341_, new_n4983_, new_n1938_, new_n169_, new_n4580_, new_n429_, new_n3927_, new_n783_, new_n1066_, v[1], new_n1744_, new_n262_, new_n5714_, new_n1263_, new_n3485_, y[2], new_n244_, new_n1504_, new_n228_, new_n1012_, new_n95_, new_n5800_, new_n493_, new_n649_, new_n121_, new_n5156_, new_n1753_, new_n3787_, new_n469_, new_n1892_, new_n257_, new_n986_, new_n133_, new_n524_, new_n82_, new_n4559_, new_n1568_, new_n3480_, new_n1649_, new_n3320_, new_n363_, new_n723_, new_n338_, new_n813_, new_n378_, new_n1678_, new_n150_, new_n937_, new_n481_, new_n3544_, new_n382_, new_n3255_, new_n381_, new_n1963_, new_n1225_, new_n1551_, new_n1047_, new_n4506_, new_n395_, new_n1835_, new_n1337_, new_n2992_, new_n207_, new_n2799_, new_n389_, new_n1046_, new_n142_, new_n5030_, new_n151_, new_n4802_, new_n267_, new_n1607_, new_n118_, new_n725_, new_n154_, new_n308_, new_n250_, new_n809_, new_n1580_, new_n1848_, new_n86_, new_n4253_, new_n796_, new_n1406_, new_n85_, new_n353_, new_n1620_, new_n127_, new_n5422_, new_n371_, new_n5069_, new_n578_, new_n4353_, new_n744_, new_n1964_, new_n953_, new_n2617_, new_n1181_, new_n1583_, new_n321_, new_n2796_, new_n137_, new_n1910_, new_n178_, new_n1825_, new_n168_, new_n5818_, new_n4584_, new_n407_, new_n3617_, new_n342_, new_n2110_, new_n230_, new_n5745_, new_n805_, new_n6087_, new_n278_, new_n593_, new_n6220_, new_n1183_, new_n1738_, new_n218_, new_n1043_, new_n140_, new_n1564_, new_n1033_, new_n1231_, new_n2908_, new_n626_, new_n1810_, new_n174_, new_n5862_, new_n161_, new_n5622_, new_n285_, new_n762_, new_n101_, new_n445_, new_n1029_, new_n313_, new_n1152_, new_n2905_, new_n208_, new_n1226_, new_n183_, new_n5074_, new_n237_, new_n311_, new_n134_, new_n4959_, new_n269_, new_n571_, new_n84_, new_n4407_, new_n83_, new_n1437_, new_n530_, new_n4249_, new_n760_, new_n3062_, new_n695_, new_n739_, new_n179_, new_n5797_, new_n2365_, new_n131_, new_n3043_, new_n171_, new_n5505_, new_n258_, new_n909_, new_n5928_, new_n164_, new_n4066_, new_n2441_, new_n369_, new_n2706_, new_n6234_, new_n270_, new_n1911_, new_n344_, new_n5371_, new_n557_, new_n752_, new_n1072_, new_n3308_, new_n459_, new_n2158_, new_n260_, new_n5481_, new_n409_, new_n4530_, new_n190_, new_n4657_, new_n523_, new_n5362_, new_n295_, new_n359_, new_n500_, new_n1922_, new_n116_, new_n753_, new_n189_, new_n6105_, new_n223_, new_n4742_, new_n255_, new_n5508_, new_n651_, new_n2497_, new_n214_, new_n1209_, new_n170_, new_n1336_, new_n275_, new_n4881_, new_n635_, new_n1166_, new_n265_, new_n365_, new_n305_, new_n2849_, new_n1258_, new_n5005_, x[1], new_n284_, new_n972_, new_n713_, new_n1700_, new_n943_, new_n5594_, new_n79_, new_n2801_, new_n239_, new_n4542_, new_n312_, new_n747_, new_n191_, new_n202_, new_n316_, new_n2804_, new_n414_, new_n1087_, new_n1165_, new_n2425_, new_n350_, new_n4481_, new_n496_, new_n4951_, new_n501_, new_n612_, new_n536_, new_n4445_, new_n355_, new_n5414_, new_n96_, new_n2473_, new_n159_, new_n836_, new_n155_, new_n1116_, new_n673_, new_n3753_, new_n128_, new_n4468_, new_n448_, new_n722_, new_n184_, new_n5918_, new_n123_, new_n5743_, new_n213_, new_n2817_, new_n268_, new_n1074_, new_n90_, new_n758_, new_n3603_, new_n6225_, new_n167_, new_n1411_, new_n87_, new_n300_, new_n560_, new_n450_, new_n1820_, new_n263_, new_n3201_, new_n157_, new_n5793_, new_n241_, new_n2705_, new_n173_, new_n5988_, new_n602_, new_n1898_, new_n334_, new_n2754_, new_n246_, new_n4508_, new_n280_, new_n1850_, new_n503_, new_n621_, new_n196_, new_n5346_, new_n144_, new_n3080_, new_n194_, new_n201_, new_n217_, new_n336_, new_n529_, new_n182_, new_n1747_, new_n346_, new_n1499_, new_n6252_, new_n129_, new_n3207_, new_n187_, new_n1584_, new_n2812_, new_n115_, new_n5158_, new_n438_, new_n5938_, new_n1135_, new_n3789_, new_n254_, new_n617_, new_n2369_, new_n238_, new_n5569_, new_n175_, new_n2749_})
361'b11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????0?????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????0???????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[3] = 1'b1;
361'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????? : coef[3] = 1'b1;
361'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????? : coef[3] = 1'b1;
361'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? : coef[3] = 1'b1;
361'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[3] = 1'b1;
361'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[3] = 1'b1;
default : coef[3] = 1'b0;
endcase
casez ({new_n525_, new_n1622_, new_n176_, new_n3741_, new_n220_, new_n3626_, new_n177_, new_n597_, new_n796_, new_n267_, new_n4374_, new_n286_, new_n5177_, new_n225_, new_n5650_, new_n221_, new_n1572_, new_n1804_, new_n2143_, new_n265_, new_n416_, new_n244_, new_n4265_, new_n360_, new_n3295_, new_n194_, new_n2708_, new_n131_, new_n4096_, new_n1889_, new_n1963_, new_n868_, new_n2582_, new_n1057_, new_n2916_, new_n341_, new_n546_, new_n6049_, new_n81_, new_n758_, y[0], new_n3762_, new_n97_, new_n3652_, new_n486_, new_n756_, new_n185_, new_n2522_, new_n487_, new_n4673_, new_n1523_, new_n277_, new_n821_, new_n472_, new_n1808_, new_n440_, new_n4574_, new_n4600_, new_n556_, new_n979_, new_n494_, new_n632_, new_n950_, new_n3378_, new_n191_, new_n1272_, new_n405_, new_n4139_, new_n671_, new_n3357_, new_n162_, new_n2564_, new_n6253_, new_n447_, new_n4213_, new_n473_, new_n742_, new_n744_, new_n1385_, new_n553_, new_n2988_, new_n605_, new_n1651_, new_n537_, new_n4444_, new_n262_, new_n5738_, u[1], new_n1001_, new_n1171_, new_n127_, new_n5149_, new_n388_, new_n2843_, new_n150_, new_n2668_, new_n469_, new_n611_, new_n442_, new_n3322_, new_n988_, new_n3147_, new_n493_, new_n3392_, new_n317_, new_n735_, new_n228_, new_n5053_, new_n299_, new_n3403_, new_n856_, new_n3673_, new_n786_, new_n3521_, new_n86_, new_n338_, new_n371_, new_n118_, new_n1431_, new_n321_, new_n5061_, new_n404_, new_n495_, new_n238_, new_n4336_, new_n578_, new_n4209_, new_n776_, new_n2839_, new_n551_, new_n5703_, new_n391_, new_n855_, new_n2275_, new_n104_, new_n4945_, new_n166_, new_n5143_, x[1], new_n230_, new_n462_, new_n1349_, new_n2926_, new_n218_, new_n4003_, new_n418_, new_n2153_, new_n132_, new_n4516_, new_n106_, new_n435_, new_n85_, new_n5667_, new_n179_, new_n1515_, new_n2420_, new_n1454_, new_n2159_, new_n171_, new_n5532_, new_n523_, new_n1508_, new_n2901_, new_n1059_, new_n2936_, new_n2896_, new_n934_, new_n1825_, new_n161_, new_n4703_, new_n311_, new_n4289_, new_n234_, new_n4651_, new_n427_, new_n2222_, new_n445_, new_n544_, new_n313_, new_n520_, new_n2567_, new_n6217_, new_n184_, new_n5726_, new_n229_, new_n1226_, new_n200_, new_n6070_, new_n306_, new_n1145_, new_n164_, new_n5947_, new_n168_, new_n5524_, new_n956_, new_n1002_, new_n196_, new_n2605_, new_n5437_, new_n336_, new_n5731_, new_n530_, new_n688_, new_n393_, new_n1722_, new_n266_, new_n1468_, new_n324_, new_n3087_, new_n140_, new_n5415_, new_n151_, new_n5072_, new_n237_, new_n1925_, new_n89_, new_n4234_, new_n183_, new_n831_, new_n187_, new_n4762_, new_n224_, new_n5739_, new_n683_, new_n1911_, new_n1463_, new_n2939_, new_n281_, new_n1007_, new_n169_, new_n3058_, new_n152_, new_n3732_, new_n92_, new_n103_, new_n303_, new_n129_, new_n718_, new_n417_, new_n5207_, new_n497_, new_n3569_, new_n157_, new_n5630_, new_n160_, new_n5602_, new_n242_, new_n5858_, new_n923_, new_n1592_, new_n272_, new_n1546_, new_n6174_, new_n173_, new_n5464_, new_n158_, new_n586_, new_n1019_, new_n1636_, new_n202_, new_n1893_, new_n397_, new_n2716_, new_n635_, new_n673_, new_n90_, new_n1481_, new_n190_, new_n5776_, new_n532_, new_n3118_, new_n189_, new_n5333_, v[0], new_n1444_, new_n438_, new_n2254_, new_n253_, new_n1998_, new_n355_, new_n448_, u[2], new_n232_, new_n2526_, new_n159_, new_n702_, new_n259_, new_n4420_, new_n296_, new_n322_, new_n315_, new_n946_, new_n365_, new_n4903_, new_n419_, new_n3014_, new_n239_, new_n1008_, new_n384_, new_n3293_, new_n155_, new_n6102_, new_n149_, new_n5744_, u[0], new_n3679_, new_n174_, new_n6167_, new_n120_, new_n2805_, new_n289_, new_n5668_, new_n385_, new_n6090_, new_n144_, new_n4055_, new_n2885_, new_n529_, new_n602_, new_n145_, new_n5657_, new_n334_, new_n612_, new_n208_, new_n5684_, new_n424_, new_n4825_, new_n554_, new_n2836_, new_n188_, new_n4957_, new_n198_, new_n3249_, new_n457_, new_n3583_, new_n318_, new_n3190_, new_n479_, new_n1040_, new_n167_, new_n4824_, new_n245_, new_n251_, new_n344_, new_n5910_, new_n254_, new_n1328_, new_n209_, new_n1714_, new_n175_, new_n3321_, new_n293_, new_n470_, new_n115_, new_n5868_, new_n2369_, new_n347_, new_n1074_, new_n697_, new_n1110_, new_n214_, new_n2135_, new_n275_, new_n5219_, new_n199_, new_n4844_})
366'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????0?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110?????????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[4] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????? : coef[4] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[4] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[4] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[4] = 1'b0;
default : coef[4] = 1'b1;
endcase
casez ({new_n1030_, new_n1267_, new_n584_, new_n1170_, new_n1195_, new_n1631_, new_n166_, new_n3217_, new_n176_, new_n2336_, new_n480_, new_n3047_, new_n1429_, new_n3587_, new_n360_, new_n2649_, new_n262_, new_n1352_, new_n122_, new_n1048_, new_n225_, new_n5829_, new_n899_, new_n1821_, new_n220_, new_n5100_, new_n1022_, new_n4284_, new_n522_, new_n1371_, new_n247_, new_n2702_, new_n228_, new_n2578_, new_n789_, new_n4305_, new_n207_, new_n5208_, new_n195_, new_n5831_, new_n748_, new_n4224_, new_n244_, new_n1806_, new_n299_, new_n1462_, v[1], new_n283_, new_n2913_, new_n498_, new_n3435_, new_n2314_, new_n1013_, new_n1175_, new_n486_, new_n5521_, new_n277_, new_n2522_, new_n94_, new_n699_, new_n387_, new_n1107_, y[0], new_n118_, new_n542_, new_n437_, new_n2648_, new_n971_, new_n1881_, new_n139_, new_n421_, new_n191_, new_n3599_, new_n2461_, new_n504_, new_n1622_, new_n403_, new_n1928_, new_n241_, new_n3993_, new_n441_, new_n1959_, new_n321_, new_n908_, new_n356_, new_n1716_, new_n454_, new_n5028_, new_n447_, new_n3117_, new_n371_, new_n742_, new_n719_, new_n2792_, new_n377_, new_n1179_, new_n353_, new_n1651_, new_n605_, new_n2584_, new_n271_, new_n4442_, new_n330_, new_n1160_, new_n578_, new_n1172_, new_n151_, new_n5081_, new_n1704_, new_n2762_, new_n725_, new_n783_, new_n339_, new_n581_, new_n465_, new_n988_, new_n524_, new_n1173_, new_n417_, new_n2787_, new_n398_, new_n1471_, new_n517_, new_n987_, new_n212_, new_n3678_, new_n148_, new_n4458_, new_n875_, new_n2742_, new_n267_, new_n3403_, new_n392_, new_n5171_, new_n459_, new_n460_, y[1], new_n4975_, new_n493_, new_n1729_, new_n619_, new_n2138_, new_n405_, new_n582_, new_n796_, new_n3554_, new_n257_, new_n2794_, new_n209_, new_n4626_, new_n86_, new_n5033_, new_n5451_, new_n154_, new_n4744_, new_n281_, new_n5916_, new_n551_, new_n565_, new_n1702_, new_n3326_, new_n226_, new_n1833_, new_n462_, new_n4310_, new_n379_, new_n4894_, new_n284_, new_n5150_, new_n413_, new_n5840_, new_n242_, new_n6125_, new_n943_, new_n1525_, new_n177_, new_n5515_, v[0], new_n2596_, new_n223_, new_n6083_, new_n203_, new_n1373_, new_n84_, new_n3754_, new_n265_, new_n1503_, new_n6277_, new_n159_, new_n1628_, new_n5922_, new_n386_, new_n666_, new_n261_, new_n664_, new_n989_, new_n3547_, new_n767_, new_n3213_, new_n279_, new_n901_, new_n342_, new_n2118_, new_n1198_, new_n184_, new_n468_, u[2], new_n1721_, new_n235_, new_n4553_, new_n270_, new_n4874_, new_n269_, new_n3612_, new_n5928_, new_n1102_, new_n5093_, new_n775_, new_n3227_, new_n1020_, new_n3985_, new_n491_, new_n5109_, new_n1137_, new_n3606_, new_n162_, new_n5966_, new_n88_, new_n5623_, new_n168_, new_n2749_, new_n249_, new_n3907_, new_n167_, new_n4154_, new_n140_, new_n5617_, new_n313_, new_n1866_, new_n172_, new_n4298_, new_n204_, new_n1105_, new_n218_, new_n5583_, new_n224_, new_n580_, new_n295_, new_n990_, new_n376_, new_n708_, new_n383_, new_n1343_, new_n427_, new_n2669_, new_n254_, new_n514_, new_n152_, new_n5166_, new_n144_, new_n5477_, new_n263_, new_n5015_, new_n557_, new_n2920_, new_n278_, new_n4806_, new_n104_, new_n981_, new_n103_, new_n5251_, new_n502_, new_n1542_, new_n98_, new_n1890_, new_n205_, new_n4960_, new_n240_, new_n1466_, new_n230_, new_n4845_, new_n155_, new_n740_, new_n727_, new_n3280_, new_n2193_, new_n6174_, new_n274_, new_n4999_, new_n287_, new_n4671_, new_n6261_, new_n173_, new_n5854_, new_n286_, new_n5814_, new_n236_, new_n4428_, new_n635_, new_n4251_, new_n129_, new_n2675_, new_n801_, new_n3688_, new_n401_, new_n5674_, new_n490_, new_n1186_, new_n161_, new_n5808_, new_n259_, new_n675_, new_n1097_, new_n3093_, new_n123_, new_n5460_, new_n256_, new_n4853_, new_n210_, new_n3323_, new_n6162_, new_n598_, new_n4849_, new_n520_, new_n2997_, new_n532_, new_n4667_, new_n1054_, new_n1815_, new_n83_, new_n276_, new_n364_, new_n190_, new_n215_, new_n411_, new_n325_, new_n872_, new_n198_, new_n1475_, new_n1575_, new_n4451_, new_n2437_, new_n229_, new_n1834_, new_n380_, new_n1501_, new_n300_, new_n1584_, new_n89_, new_n2830_, new_n200_, new_n5182_, new_n6270_, new_n355_, new_n1362_, new_n326_, new_n2520_, new_n1986_, new_n201_, new_n4136_, new_n753_, new_n2126_, new_n79_, new_n672_, new_n1095_, new_n1919_, new_n3067_, new_n2063_, new_n1561_, new_n3260_, new_n183_, new_n5601_, new_n2888_, new_n246_, new_n851_, new_n1348_, new_n3138_, new_n479_, new_n906_, new_n993_, new_n6077_, new_n157_, new_n5398_, new_n531_, new_n1714_, new_n199_, new_n2679_})
387'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????011?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????? : coef[5] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????? : coef[5] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00?????? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???? : coef[5] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[5] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[5] = 1'b0;
default : coef[5] = 1'b1;
endcase
casez ({new_n101_, new_n220_, new_n3597_, new_n127_, new_n5244_, new_n299_, new_n1138_, new_n6268_, new_n2513_, new_n3627_, new_n262_, new_n2261_, new_n305_, new_n1242_, new_n1886_, new_n4020_, new_n306_, new_n4438_, new_n140_, new_n1596_, new_n171_, new_n2711_, new_n177_, new_n374_, new_n223_, new_n6008_, new_n270_, new_n770_, new_n86_, new_n2429_, new_n168_, new_n4562_, new_n250_, new_n724_, new_n342_, new_n4915_, new_n484_, new_n797_, new_n170_, new_n577_, new_n153_, new_n5203_, new_n112_, new_n1877_, new_n311_, new_n1177_, new_n284_, new_n5784_, new_n438_, new_n2818_, new_n239_, new_n5483_, new_n584_, new_n3569_, new_n6258_, new_n83_, new_n3838_, new_n781_, new_n3192_, new_n242_, new_n1411_, new_n636_, new_n2969_, new_n432_, new_n3029_, new_n166_, new_n5798_, new_n188_, new_n4465_, new_n2890_, new_n176_, new_n1569_, new_n173_, new_n5155_, new_n160_, new_n2646_, new_n103_, new_n2115_, new_n230_, new_n1718_, new_n175_, new_n3638_, new_n190_, new_n2627_, new_n186_, new_n1352_, new_n623_, new_n1396_, new_n198_, new_n2657_, new_n326_, new_n1885_, new_n158_, new_n5395_, new_n90_, new_n1672_, new_n236_, new_n673_, new_n162_, new_n1209_, new_n123_, new_n5546_, new_n2479_, new_n267_, new_n477_, new_n634_, new_n1388_, new_n632_, new_n1956_, new_n225_, new_n2299_, new_n766_, new_n938_, new_n82_, new_n699_, new_n865_, new_n3234_, new_n2324_, new_n241_, new_n908_, new_n214_, new_n1713_, new_n976_, new_n3104_, new_n486_, new_n4614_, new_n671_, new_n1338_, new_n191_, new_n826_, new_n958_, new_n3557_, new_n248_, new_n3826_, new_n4647_, new_n555_, new_n1639_, new_n121_, new_n2664_, new_n142_, new_n1202_, new_n164_, new_n1022_, new_n179_, new_n5899_, new_n210_, new_n760_, new_n161_, new_n4804_, new_n370_, new_n468_, new_n1237_, new_n463_, new_n3208_, new_n132_, new_n506_, new_n6216_, new_n6255_, new_n232_, new_n3103_, new_n557_, new_n3140_, new_n155_, new_n1564_, new_n255_, new_n1530_, new_n240_, new_n5312_, new_n608_, new_n1019_, new_n216_, new_n3430_, new_n318_, new_n4768_, new_n682_, new_n2512_, new_n448_, new_n697_, new_n791_, new_n1640_, new_n144_, new_n1806_, new_n234_, new_n4865_, new_n185_, new_n2599_, new_n205_, new_n5367_, new_n471_, new_n3010_, new_n598_, new_n1523_, new_n145_, new_n6110_, new_n277_, new_n4554_, new_n1276_, new_n1606_, new_n189_, new_n3240_, new_n556_, new_n3946_, new_n515_, new_n1932_, new_n184_, new_n2775_, new_n1353_, new_n1539_, new_n361_, new_n3711_, new_n334_, new_n442_, new_n319_, new_n4328_, new_n389_, new_n868_, new_n271_, new_n1952_, new_n605_, new_n3691_, new_n786_, new_n3022_, new_n366_, new_n5038_, new_n371_, new_n957_, new_n377_, new_n1635_, new_n1867_, new_n1961_, new_n196_, new_n1755_, new_n430_, new_n1062_, new_n309_, new_n5236_, new_n725_, new_n1804_, new_n417_, new_n1211_, new_n606_, new_n2756_, new_n247_, new_n1108_, new_n317_, new_n2117_, new_n1035_, new_n3577_, new_n541_, new_n1067_, new_n154_, new_n5183_, new_n115_, new_n1723_, new_n405_, new_n4230_, new_n118_, new_n1472_, new_n85_, new_n5187_, new_n169_, new_n204_, new_n437_, new_n360_, new_n1839_, new_n1726_, new_n2912_, new_n6188_, new_n719_, new_n1717_, new_n139_, new_n4627_, new_n295_, new_n744_, new_n5675_, new_n460_, new_n2732_, new_n749_, new_n1871_, new_n3320_, new_n3581_, new_n307_, new_n3962_, new_n393_, new_n1903_, new_n266_, new_n4028_, new_n456_, new_n1366_, new_n919_, new_n368_, new_n3848_, new_n113_, new_n5516_, new_n89_, new_n866_, new_n424_, new_n1983_, new_n167_, new_n1786_, new_n172_, new_n4056_, new_n151_, new_n3370_, new_n1200_, new_n1813_, new_n709_, new_n1503_, new_n683_, new_n869_, new_n346_, new_n642_, new_n1040_, new_n2838_, new_n238_, new_n375_, new_n84_, new_n4897_, new_n187_, new_n643_, new_n253_, new_n1326_, new_n315_, new_n5366_, new_n245_, new_n603_, new_n336_, new_n6103_, new_n296_, new_n5185_, new_n251_, new_n289_, new_n511_, new_n1015_, new_n679_, new_n1161_, v[2], new_n4185_, new_n1794_, new_n6290_, new_n6246_, new_n6269_})
342'b011??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[6] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? : coef[6] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?? : coef[6] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0? : coef[6] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0 : coef[6] = 1'b1;
default : coef[6] = 1'b0;
endcase
casez ({new_n278_, new_n6107_, new_n247_, new_n2594_, new_n221_, new_n2619_, new_n127_, new_n4068_, new_n267_, new_n6079_, new_n121_, new_n4953_, new_n265_, new_n3548_, new_n829_, new_n1487_, new_n1138_, new_n1812_, new_n597_, new_n4604_, new_n220_, new_n5530_, new_n161_, new_n3836_, new_n742_, new_n864_, new_n748_, new_n1948_, new_n192_, new_n5137_, new_n1119_, new_n2927_, new_n135_, new_n2146_, new_n522_, new_n2556_, new_n98_, new_n292_, new_n2551_, new_n698_, new_n1093_, new_n345_, new_n387_, new_n122_, new_n911_, new_n228_, new_n5029_, new_n486_, new_n1254_, new_n331_, new_n2676_, new_n1029_, new_n1338_, new_n1152_, v[2], new_n2586_, new_n360_, new_n1456_, u[0], new_n4335_, new_n5434_, new_n1434_, new_n225_, new_n3675_, new_n219_, new_n5771_, new_n276_, new_n807_, new_n215_, new_n668_, new_n1148_, new_n3098_, new_n96_, new_n3933_, new_n248_, new_n4338_, new_n1188_, new_n82_, new_n879_, new_n101_, new_n3807_, new_n290_, new_n4387_, new_n776_, new_n868_, new_n606_, new_n3105_, new_n371_, new_n4475_, new_n980_, new_n2928_, new_n358_, new_n1483_, new_n214_, new_n2793_, new_n183_, new_n1357_, new_n783_, new_n1725_, new_n430_, new_n904_, new_n388_, new_n809_, new_n216_, new_n1063_, new_n1288_, new_n329_, new_n1883_, new_n508_, new_n1150_, new_n1236_, new_n2171_, new_n622_, new_n1001_, new_n1065_, new_n3197_, new_n633_, new_n2768_, new_n6254_, new_n459_, new_n744_, u[1], new_n309_, new_n953_, new_n578_, new_n1557_, new_n2367_, new_n711_, new_n3264_, new_n712_, new_n2829_, new_n537_, new_n3759_, new_n579_, new_n1073_, new_n447_, new_n3863_, new_n356_, new_n3818_, new_n6236_, new_n616_, new_n5833_, new_n1646_, new_n1941_, new_n391_, new_n3450_, new_n284_, new_n643_, new_n103_, new_n2674_, new_n164_, new_n4770_, new_n306_, new_n2061_, new_n565_, new_n2941_, new_n230_, new_n1731_, new_n226_, new_n5913_, new_n137_, new_n5326_, new_n104_, new_n5856_, new_n166_, new_n6026_, new_n176_, new_n5510_, new_n218_, new_n5565_, new_n242_, new_n6089_, new_n618_, new_n4397_, new_n5927_, new_n150_, new_n2834_, new_n2904_, new_n132_, new_n1203_, new_n134_, new_n644_, new_n179_, new_n2110_, new_n171_, new_n1481_, new_n279_, new_n1112_, new_n223_, new_n5643_, new_n484_, new_n3492_, new_n2406_, new_n269_, new_n5607_, new_n501_, new_n1403_, new_n311_, new_n3873_, new_n368_, new_n1163_, new_n172_, new_n947_, new_n448_, new_n5377_, new_n113_, new_n3474_, new_n210_, new_n915_, new_n1373_, new_n1640_, new_n369_, new_n1907_, new_n283_, new_n3471_, new_n342_, new_n2222_, new_n393_, new_n5249_, new_n231_, new_n2565_, new_n266_, new_n419_, new_n307_, new_n3806_, new_n191_, new_n775_, new_n504_, new_n800_, new_n140_, new_n5276_, new_n208_, new_n710_, new_n385_, new_n2429_, new_n1174_, new_n3179_, new_n1567_, new_n2777_, new_n300_, new_n1556_, new_n168_, new_n5806_, new_n6267_, new_n237_, new_n446_, new_n313_, new_n5908_, new_n427_, new_n1348_, new_n527_, new_n990_, new_n285_, new_n2577_, new_n375_, new_n1110_, new_n732_, new_n794_, new_n118_, new_n5656_, new_n272_, new_n5740_, new_n551_, new_n701_, new_n3881_, new_n239_, new_n3068_, new_n409_, new_n964_, new_n155_, new_n804_, new_n289_, new_n2502_, new_n145_, new_n5642_, new_n232_, new_n734_, new_n871_, new_n1176_, new_n157_, new_n891_, new_n529_, new_n1543_, new_n500_, new_n2055_, new_n438_, new_n1627_, new_n2570_, new_n418_, new_n1381_, new_n160_, new_n5917_, new_n287_, new_n2574_, new_n209_, new_n1209_, new_n123_, new_n5107_, new_n2193_, new_n249_, new_n1485_, new_n509_, new_n1210_, new_n467_, new_n1016_, new_n178_, new_n5164_, new_n158_, new_n4469_, new_n236_, new_n1733_, new_n280_, new_n4477_, new_n170_, new_n895_, new_n159_, new_n2993_, new_n188_, new_n414_, new_n682_, new_n1379_, new_n175_, new_n5597_, new_n433_, new_n3045_, new_n303_, new_n1642_, new_n917_, new_n3030_, new_n478_, new_n5525_, new_n255_, new_n544_, new_n318_, new_n2127_, new_n496_, new_n672_, new_n186_, new_n3426_, new_n650_, new_n955_, new_n426_, new_n962_, new_n84_, new_n4606_, new_n174_, new_n6200_, new_n2853_, new_n355_, new_n454_, new_n602_, new_n1135_, new_n245_, new_n1699_, new_n336_, new_n722_, new_n323_, new_n5606_, new_n88_, new_n4641_, new_n189_, new_n4320_, new_n324_, new_n2399_, new_n167_, new_n6086_, new_n263_, new_n5495_, new_n291_, new_n3139_, new_n1305_, new_n3404_, new_n204_, new_n1747_, new_n363_, new_n2788_, new_n217_, new_n862_, new_n359_, new_n2694_, new_n233_, new_n3590_, new_n673_, new_n1619_, new_n211_, new_n1458_, new_n187_, new_n4112_, new_n254_, new_n5394_, new_n205_, new_n3994_})
392'b10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????110????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????1??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????1????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????0??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????? : coef[7] = 1'b0;
392'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????? : coef[7] = 1'b0;
392'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???? : coef[7] = 1'b0;
392'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[7] = 1'b0;
392'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[7] = 1'b0;
default : coef[7] = 1'b1;
endcase
casez ({new_n166_, new_n988_, new_n221_, new_n1026_, new_n286_, new_n3905_, new_n225_, new_n5999_, new_n267_, new_n5159_, new_n82_, new_n1520_, new_n384_, new_n3241_, new_n2040_, new_n699_, new_n2505_, new_n121_, new_n614_, new_n262_, new_n4747_, new_n4600_, new_n220_, new_n1502_, new_n169_, new_n649_, new_n1600_, new_n3143_, new_n191_, new_n5099_, new_n1376_, new_n3121_, new_n874_, new_n2654_, new_n579_, new_n1881_, new_n522_, new_n5357_, new_n214_, new_n5264_, new_n148_, new_n5041_, new_n430_, new_n1154_, new_n441_, new_n1926_, new_n372_, new_n382_, new_n142_, new_n4724_, new_n94_, new_n5557_, new_n127_, new_n5528_, new_n742_, new_n1103_, new_n353_, new_n957_, new_n290_, new_n1390_, new_n2245_, new_n524_, new_n1948_, new_n381_, new_n3718_, new_n677_, new_n2517_, new_n310_, new_n987_, new_n999_, new_n1621_, new_n309_, new_n3912_, new_n821_, new_n3914_, new_n4639_, new_n95_, new_n859_, new_n6184_, new_n725_, new_n4577_, new_n150_, new_n2807_, new_n465_, new_n1030_, new_n377_, new_n1046_, new_n6279_, new_n1067_, new_n3119_, new_n395_, new_n3536_, new_n343_, new_n980_, new_n207_, new_n975_, new_n212_, new_n2796_, new_n676_, new_n2154_, new_n1723_, new_n4384_, new_n1472_, new_n1955_, u[0], new_n122_, new_n950_, new_n154_, new_n5480_, new_n327_, new_n875_, new_n1001_, new_n3461_, new_n460_, new_n3981_, new_n787_, new_n1132_, new_n371_, new_n3686_, new_n339_, new_n3702_, new_n319_, new_n1479_, new_n455_, new_n3849_, new_n423_, new_n1807_, new_n1222_, new_n2981_, new_n1583_, new_n2767_, new_n1568_, new_n2780_, new_n218_, new_n1727_, new_n137_, new_n1461_, new_n2900_, new_n230_, new_n374_, new_n168_, new_n1345_, new_n153_, new_n3061_, new_n164_, new_n5018_, new_n902_, new_n3006_, new_n2298_, new_n86_, new_n6139_, new_n6232_, new_n456_, new_n3469_, new_n642_, new_n4231_, new_n6031_, new_n644_, new_n1183_, new_n805_, new_n2164_, new_n1059_, new_n3314_, new_n171_, new_n6007_, new_n266_, new_n6063_, new_n6033_, new_n179_, new_n475_, new_n306_, new_n1915_, new_n2279_, new_n159_, new_n5459_, new_n261_, new_n5154_, new_n6208_, new_n546_, new_n2109_, new_n140_, new_n5919_, new_n285_, new_n463_, new_n313_, new_n2326_, new_n435_, new_n3162_, new_n174_, new_n4871_, new_n112_, new_n3327_, new_n461_, new_n810_, new_n215_, new_n5857_, new_n270_, new_n1168_, new_n496_, new_n5293_, new_n1545_, new_n1878_, new_n323_, new_n4421_, new_n89_, new_n1731_, new_n602_, new_n1403_, new_n1615_, new_n3271_, new_n1000_, new_n4759_, new_n334_, new_n4120_, new_n200_, new_n6106_, new_n324_, new_n3506_, new_n113_, new_n4772_, new_n2441_, new_n151_, new_n5994_, new_n503_, new_n5691_, new_n183_, new_n5826_, new_n237_, new_n3760_, new_n4638_, new_n235_, new_n3414_, new_n224_, new_n5632_, new_n530_, new_n1151_, new_n187_, new_n6073_, new_n342_, new_n5259_, new_n583_, new_n1652_, new_n260_, new_n4920_, new_n190_, new_n6003_, new_n284_, new_n4763_, new_n259_, new_n2795_, new_n239_, new_n1790_, new_n135_, new_n1399_, new_n528_, new_n4513_, new_n103_, new_n2604_, new_n194_, new_n1890_, new_n176_, new_n1448_, new_n359_, new_n646_, new_n497_, new_n1311_, new_n380_, new_n2113_, new_n242_, new_n661_, new_n205_, new_n4099_, new_n808_, new_n1814_, new_n177_, new_n5706_, new_n467_, new_n1129_, new_n420_, new_n3534_, new_n162_, new_n5215_, new_n255_, new_n1112_, new_n607_, new_n960_, v[1], new_n87_, new_n352_, new_n272_, new_n5613_, new_n170_, new_n5121_, v[0], new_n96_, new_n124_, new_n139_, new_n265_, new_n1074_, new_n2714_, new_n4610_, new_n178_, new_n6171_, new_n2479_, new_n246_, new_n5672_, new_n621_, new_n4416_, new_n161_, new_n861_, new_n297_, new_n1038_, new_n289_, new_n3286_, new_n1097_, new_n1499_, new_n354_, new_n3519_, new_n210_, new_n2753_, new_n195_, new_n202_, new_n458_, new_n729_, new_n189_, new_n5262_, new_n292_, new_n1575_, new_n123_, new_n1008_, new_n498_, new_n3423_, new_n129_, new_n185_, new_n2488_, new_n144_, new_n5825_, new_n175_, new_n5410_, new_n743_, new_n3483_, new_n268_, new_n5467_, new_n173_, new_n5883_, new_n5440_, new_n479_, new_n556_, new_n1054_, new_n2950_, new_n312_, new_n454_, new_n325_, new_n4936_, new_n410_, new_n2972_, new_n208_, new_n1056_, new_n424_, new_n1071_, new_n280_, new_n4696_, new_n88_, new_n5934_, new_n450_, new_n2068_, new_n145_, new_n5351_, new_n196_, new_n5654_, new_n355_, new_n873_, new_n346_, new_n2155_, new_n157_, new_n1274_, new_n628_, new_n2819_, new_n263_, new_n1590_, new_n704_, new_n1194_, new_n2888_, new_n318_, new_n1831_, new_n251_, new_n2555_, new_n182_, new_n4925_, new_n204_, new_n5258_, new_n274_, new_n4776_, new_n1709_, new_n2773_, new_n258_, new_n4496_, new_n1096_, new_n3655_})
399'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1011?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[8] = 1'b1;
399'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????? : coef[8] = 1'b1;
399'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???? : coef[8] = 1'b1;
399'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[8] = 1'b1;
399'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[8] = 1'b1;
default : coef[8] = 1'b0;
endcase
casez ({new_n480_, new_n5101_, new_n309_, new_n5301_, new_n351_, new_n1921_, new_n221_, new_n4644_, new_n220_, new_n2616_, new_n1869_, new_n3235_, new_n299_, new_n4746_, new_n488_, new_n2588_, new_n1711_, new_n5181_, new_n416_, new_n3580_, new_n139_, new_n678_, new_n988_, new_n2948_, new_n102_, new_n143_, new_n165_, new_n150_, new_n4306_, new_n430_, new_n4994_, new_n671_, new_n1800_, new_n388_, new_n1154_, new_n2907_, new_n6287_, new_n229_, new_n5397_, new_n1132_, new_n3727_, new_n328_, new_n1360_, new_n469_, new_n2841_, new_n454_, new_n1075_, new_n121_, new_n1615_, new_n103_, new_n432_, new_n1034_, new_n95_, new_n1866_, new_n503_, new_n1413_, new_n723_, new_n2937_, new_n249_, new_n809_, new_n295_, new_n453_, new_n94_, new_n1859_, new_n6282_, new_n335_, new_n4133_, new_n5675_, new_n435_, new_n1882_, new_n82_, new_n2825_, new_n323_, new_n2958_, new_n764_, new_n2618_, new_n225_, new_n3462_, new_n228_, new_n5428_, new_n5445_, new_n2858_, new_n6230_, new_n1035_, new_n4271_, new_n154_, new_n2793_, new_n254_, new_n816_, new_n343_, new_n953_, new_n369_, new_n2130_, new_n431_, new_n4655_, new_n524_, new_n5266_, new_n115_, new_n5673_, new_n251_, new_n2259_, new_n271_, new_n790_, new_n80_, new_n5228_, new_n489_, new_n735_, new_n606_, new_n1646_, new_n162_, new_n1201_, new_n485_, new_n1667_, new_n311_, new_n1758_, new_n391_, new_n5220_, new_n270_, new_n2091_, new_n226_, new_n5340_, x[0], new_n86_, new_n521_, new_n6228_, new_n218_, new_n5298_, new_n724_, new_n3221_, new_n1113_, new_n1577_, new_n652_, new_n713_, new_n386_, new_n1854_, new_n774_, new_n1876_, new_n178_, new_n4870_, new_n350_, new_n5493_, new_n164_, new_n2338_, new_n302_, new_n4261_, new_n5962_, new_n168_, new_n947_, new_n5457_, new_n179_, new_n1528_, new_n5920_, new_n171_, new_n6023_, new_n6233_, new_n174_, new_n626_, new_n285_, new_n2638_, new_n313_, new_n2334_, new_n2905_, new_n183_, new_n1503_, new_n172_, new_n4964_, new_n269_, new_n5375_, new_n307_, new_n2725_, new_n2297_, new_n703_, new_n739_, new_n88_, new_n6135_, new_n695_, new_n1137_, new_n860_, new_n2515_, new_n182_, new_n5135_, new_n258_, new_n784_, new_n167_, new_n1783_, new_n187_, new_n1969_, new_n676_, new_n1773_, u[2], new_n2801_, new_n607_, new_n1165_, new_n157_, new_n1534_, new_n255_, new_n798_, new_n186_, new_n4821_, new_n123_, new_n5823_, new_n359_, new_n5774_, new_n1096_, new_n2643_, new_n291_, new_n4726_, new_n278_, new_n1208_, new_n413_, new_n1747_, new_n364_, new_n5331_, new_n265_, new_n1625_, new_n315_, new_n899_, new_n240_, new_n2814_, new_n152_, new_n2771_, new_n500_, new_n1390_, new_n281_, new_n4635_, new_n230_, new_n5025_, new_n176_, new_n1924_, new_n236_, new_n5751_, new_n242_, new_n2603_, new_n1129_, new_n1405_, new_n222_, new_n5877_, new_n771_, new_n943_, new_n1257_, new_n1475_, new_n213_, new_n5077_, new_n90_, new_n4882_, new_n190_, new_n5368_, new_n215_, new_n2609_, new_n91_, new_n2736_, new_n504_, new_n3804_, new_n536_, new_n1076_, new_n2895_, new_n241_, new_n1476_, new_n714_, new_n1311_, new_n216_, new_n3236_, new_n192_, new_n985_, new_n217_, new_n4954_, new_n144_, new_n698_, new_n185_, new_n289_, new_n356_, new_n2114_, new_n612_, new_n5407_, new_n268_, new_n502_, new_n175_, new_n1533_, new_n161_, new_n1120_, new_n420_, new_n1829_, new_n528_, new_n858_, new_n272_, new_n1820_, new_n199_, new_n4911_, new_n458_, new_n5335_, new_n189_, new_n1398_, new_n239_, new_n1904_, new_n200_, new_n5788_, new_n1298_, new_n3276_, new_n129_, new_n4326_, new_n545_, new_n3361_, new_n224_, new_n1428_, new_n1491_, new_n3101_, new_n153_, new_n4980_, new_n253_, new_n1668_, new_n2933_, new_n3318_, new_n1879_, new_n2962_})
314'b10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????111??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????001?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[9] = 1'b1;
314'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[9] = 1'b1;
314'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[9] = 1'b1;
default : coef[9] = 1'b0;
endcase
casez ({new_n184_, new_n5037_, new_n95_, new_n2595_, new_n220_, new_n1278_, new_n276_, new_n2780_, new_n426_, new_n787_, new_n346_, new_n548_, new_n317_, new_n1150_, new_n250_, new_n3791_, new_n80_, new_n133_, new_n987_, new_n1023_, new_n4650_, new_n225_, new_n5683_, u[2], new_n4632_, new_n815_, new_n1132_, new_n267_, new_n1604_, new_n127_, new_n4086_, new_n719_, new_n2117_, new_n207_, new_n4937_, new_n122_, new_n6010_, new_n118_, new_n4119_, new_n1012_, new_n3152_, new_n498_, new_n3238_, new_n2514_, new_n4815_, new_n135_, new_n1494_, new_n301_, new_n553_, new_n162_, new_n723_, new_n405_, new_n3180_, new_n339_, new_n1646_, new_n796_, new_n1892_, new_n238_, new_n4470_, new_n84_, new_n1470_, new_n387_, new_n1957_, new_n1013_, new_n4334_, new_n372_, new_n435_, new_n776_, new_n5116_, new_n605_, new_n3582_, x[1], y[2], new_n1213_, new_n1370_, new_n1867_, new_n214_, new_n1732_, new_n335_, new_n1941_, new_n6248_, new_n271_, new_n874_, new_n243_, new_n3640_, new_n82_, new_n3731_, new_n299_, new_n1123_, new_n81_, new_n762_, new_n524_, new_n2700_, new_n77_, new_n329_, new_n2499_, new_n321_, new_n975_, new_n330_, new_n790_, new_n1222_, new_n2978_, new_n473_, new_n1943_, new_n218_, new_n1665_, new_n373_, new_n751_, new_n345_, new_n990_, new_n311_, new_n1133_, new_n618_, new_n1134_, new_n564_, new_n626_, new_n451_, new_n1183_, new_n164_, new_n6149_, new_n167_, new_n978_, new_n151_, new_n6170_, new_n1169_, new_n5126_, new_n489_, new_n1463_, new_n2431_, new_n1199_, new_n2968_, new_n85_, new_n101_, new_n2680_, new_n191_, new_n386_, new_n444_, new_n171_, new_n5864_, new_n100_, new_n411_, new_n421_, new_n140_, new_n5328_, new_n183_, new_n5568_, new_n179_, new_n5429_, new_n169_, new_n4787_, new_n1004_, new_n1097_, new_n89_, new_n580_, new_n168_, new_n1361_, new_n305_, new_n577_, new_n674_, new_n2159_, new_n1239_, new_n285_, new_n384_, new_n427_, new_n2318_, new_n877_, new_n1362_, new_n269_, new_n3821_, new_n203_, new_n810_, new_n2374_, new_n146_, new_n2820_, new_n375_, new_n4711_, new_n342_, new_n2797_, new_n279_, new_n899_, new_n307_, new_n2157_, new_n199_, new_n831_, new_n2455_, new_n170_, new_n5785_, new_n153_, new_n2833_, new_n695_, new_n989_, new_n132_, new_n6132_, new_n88_, new_n841_, new_n291_, new_n845_, new_n6231_, new_n103_, new_n910_, new_n2594_, new_n3689_, new_n536_, new_n2317_, new_n149_, new_n6117_, new_n145_, new_n6119_, new_n175_, new_n939_, new_n204_, new_n3345_, new_n224_, new_n1459_, new_n174_, new_n5964_, new_n482_, new_n1815_, new_n323_, new_n612_, new_n433_, new_n3421_, new_n246_, new_n3420_, new_n187_, new_n519_, v[2], new_n4141_, new_n240_, new_n824_, new_n675_, new_n1455_, new_n257_, new_n2804_, new_n186_, new_n1826_, new_n2853_, new_n254_, new_n6094_, new_n630_, new_n1312_, new_n158_, new_n5341_, new_n161_, new_n5636_, new_n90_, new_n98_, new_n283_, new_n334_, new_n1270_, new_n281_, new_n754_, new_n176_, new_n1741_, new_n230_, new_n1221_, new_n2880_, new_n927_, new_n1760_, new_n539_, new_n3768_, new_n202_, new_n1205_, new_n107_, new_n208_, new_n1769_, new_n560_, new_n1363_, new_n607_, new_n1071_, new_n2244_, new_n4923_, new_n1486_, new_n4691_, new_n229_, new_n1072_, new_n251_, new_n410_, new_n325_, new_n3997_, new_n96_, new_n4649_, new_n280_, new_n3822_, new_n333_, new_n857_, new_n265_, new_n458_, new_n399_, new_n3935_, new_n1482_, new_n3032_, new_n192_, new_n3323_, new_n155_, new_n5372_, new_n506_, new_n1801_, new_n545_, new_n3515_, new_n241_, new_n3833_, new_n964_, new_n5695_, new_n129_, new_n4529_, new_n242_, new_n3810_, new_n157_, new_n5553_, new_n142_, new_n1736_, new_n1177_, new_n1575_, new_n255_, new_n2151_, new_n178_, new_n1830_, new_n144_, new_n331_, v[1], new_n222_, new_n472_, new_n532_, new_n1089_, new_n277_, new_n502_, new_n123_, new_n5332_, new_n190_, new_n3391_, new_n213_, new_n5610_})
333'b10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????011?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????001??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????010??????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[10] = 1'b1;
333'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[10] = 1'b1;
333'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011?????????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???? : coef[10] = 1'b1;
333'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[10] = 1'b1;
333'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[10] = 1'b1;
default : coef[10] = 1'b0;
endcase
casez ({new_n360_, new_n3310_, new_n127_, new_n2572_, new_n242_, new_n3878_, new_n548_, new_n3178_, new_n265_, new_n979_, new_n620_, new_n3786_, new_n86_, new_n978_, new_n580_, new_n1267_, new_n674_, new_n3653_, new_n379_, new_n1705_, new_n552_, new_n565_, new_n2494_, new_n1253_, new_n241_, new_n3075_, new_n168_, new_n5836_, new_n137_, new_n5108_, new_n166_, new_n6104_, new_n160_, new_n1306_, new_n153_, new_n4727_, new_n261_, new_n1118_, new_n446_, new_n3489_, new_n5659_, new_n164_, new_n5570_, new_n179_, new_n948_, new_n171_, new_n5289_, new_n783_, new_n2833_, new_n106_, new_n170_, new_n430_, new_n1578_, new_n3736_, new_n281_, new_n2830_, new_n291_, new_n584_, new_n926_, new_n1055_, new_n284_, new_n5596_, new_n232_, new_n1092_, new_n1589_, new_n2102_, new_n240_, new_n1345_, new_n464_, new_n1816_, new_n176_, new_n5404_, new_n230_, new_n5269_, new_n213_, new_n4169_, new_n2570_, new_n394_, new_n3350_, new_n528_, new_n726_, new_n129_, new_n1026_, new_n792_, new_n1129_, new_n177_, new_n5338_, new_n280_, new_n943_, new_n190_, new_n1854_, new_n6239_, new_n263_, new_n2337_, new_n1120_, new_n1540_, new_n118_, new_n1282_, new_n352_, new_n3020_, new_n444_, new_n2574_, new_n467_, new_n1162_, new_n217_, new_n1505_, new_n1210_, new_n3048_, new_n425_, new_n3250_, new_n158_, new_n811_, new_n941_, new_n3113_, new_n1485_, new_n3187_, new_n746_, new_n3191_, new_n636_, new_n805_, new_n1931_, new_n3434_, new_n397_, new_n3601_, new_n823_, new_n1709_, new_n178_, new_n595_, new_n96_, new_n3808_, new_n139_, new_n3136_, new_n210_, new_n816_, new_n767_, new_n1551_, new_n262_, new_n901_, new_n225_, new_n2302_, new_n83_, new_n4609_, new_n84_, new_n4682_, new_n6210_, new_n6259_, new_n1602_, new_n2518_, new_n442_, new_n461_, new_n247_, new_n4032_, new_n441_, new_n2677_, new_n215_, new_n1374_, new_n340_, new_n864_, new_n6032_, new_n267_, new_n1735_, new_n219_, new_n4979_, new_n249_, new_n1202_, new_n1959_, new_n5846_, new_n429_, new_n4258_, new_n122_, new_n4370_, new_n211_, new_n248_, new_n319_, new_n148_, new_n1066_, new_n226_, new_n5497_, new_n536_, new_n4893_, new_n456_, new_n682_, new_n6277_, new_n714_, new_n1158_, new_n6185_, new_n530_, new_n1915_, new_n231_, new_n4095_, new_n159_, new_n4386_, new_n1527_, new_n342_, new_n4277_, new_n307_, new_n520_, new_n172_, new_n562_, new_n279_, new_n5722_, new_n269_, new_n5682_, new_n260_, new_n1721_, new_n246_, new_n5841_, new_n161_, new_n1438_, new_n302_, new_n2683_, new_n256_, new_n490_, new_n396_, new_n1708_, new_n192_, new_n5390_, new_n5958_, new_n367_, new_n433_, new_n2488_, new_n144_, new_n6020_, new_n184_, new_n1140_, new_n205_, new_n5373_, new_n149_, new_n1399_, new_n751_, new_n4357_, new_n174_, new_n861_, new_n245_, new_n1423_, new_n259_, new_n4695_, new_n1168_, new_n2166_, new_n350_, new_n1680_, new_n3937_, new_n454_, new_n1170_, new_n275_, new_n3792_, new_n290_, new_n1634_, new_n152_, new_n1494_, new_n524_, new_n3681_, new_n324_, new_n4786_, new_n282_, new_n381_, new_n957_, new_n1703_, new_n220_, new_n1108_, new_n1061_, new_n4314_, new_n309_, new_n813_, new_n81_, new_n4739_, new_n495_, new_n1046_, new_n447_, new_n1964_, new_n142_, new_n5711_, new_n154_, new_n5815_, new_n980_, new_n1554_, new_n389_, new_n4450_, new_n162_, new_n4709_, new_n395_, new_n1639_, new_n473_, new_n5223_, new_n541_, new_n1064_, new_n243_, new_n2309_, new_n2855_, new_n299_, new_n2573_, new_n437_, new_n2131_, new_n749_, new_n2743_, new_n228_, new_n5541_, new_n187_, new_n1755_, new_n383_, new_n1073_, new_n150_, new_n5902_, new_n169_, new_n867_, new_n141_, new_n654_, new_n2529_, new_n604_, new_n1380_, new_n274_, new_n2794_, new_n77_, new_n5435_, new_n271_, new_n3984_, new_n953_, new_n2593_, new_n505_, new_n2767_, new_n1382_, new_n4455_, new_n424_, new_n618_, new_n218_, new_n5564_, new_n285_, new_n2822_, new_n131_, new_n4752_, new_n140_, new_n4205_, new_n306_, new_n5035_, new_n647_, new_n3643_, new_n201_, new_n5268_, new_n207_, new_n2706_, new_n2187_, new_n465_, new_n844_, new_n216_, new_n4563_, new_n266_, new_n1617_, new_n224_, new_n6113_, new_n132_, new_n824_, new_n391_, new_n582_, new_n270_, new_n3511_, new_n202_, new_n323_, new_n704_, new_n968_, new_n782_, new_n1541_, new_n89_, new_n5163_, new_n697_, new_n739_, new_n173_, new_n6060_, new_n200_, new_n4491_, new_n155_, new_n2623_, new_n334_, new_n4908_, new_n812_, new_n1363_, new_n189_, new_n1916_, new_n533_, new_n603_, new_n255_, new_n1847_, new_n336_, new_n5550_, new_n157_, new_n1616_, new_n167_, new_n985_, new_n151_, new_n754_, new_n503_, new_n4855_, new_n183_, new_n5951_, new_n906_, new_n1387_, new_n289_, new_n679_, new_n239_, new_n2133_, new_n251_, new_n2655_, new_n1569_, new_n3007_, new_n145_, new_n862_, new_n272_, new_n5765_, new_n175_, new_n3437_, new_n392_, new_n637_, new_n123_, new_n3901_, new_n199_, new_n623_, new_n258_, new_n2770_})
417'b11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????1???????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[11] = 1'b0;
417'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[11] = 1'b0;
417'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[11] = 1'b0;
default : coef[11] = 1'b1;
endcase
casez ({new_n103_, new_n274_, new_n480_, new_n418_, new_n1357_, new_n2211_, new_n360_, new_n3376_, new_n247_, new_n1929_, new_n228_, new_n3336_, new_n398_, new_n2758_, new_n597_, new_n4069_, new_n122_, new_n4969_, new_n5436_, new_n160_, new_n6091_, new_n168_, new_n1857_, new_n1649_, new_n4507_, new_n311_, new_n5213_, new_n734_, new_n2777_, new_n140_, new_n5662_, new_n171_, new_n1663_, new_n530_, new_n857_, new_n261_, new_n965_, new_n166_, new_n6012_, new_n2313_, new_n279_, new_n4789_, new_n391_, new_n2506_, new_n2900_, new_n409_, new_n551_, new_n131_, new_n2608_, new_n792_, new_n3477_, new_n176_, new_n2651_, new_n190_, new_n6076_, new_n202_, new_n855_, new_n144_, new_n1886_, new_n249_, new_n4755_, new_n178_, new_n5995_, new_n1019_, new_n1542_, new_n86_, new_n1555_, new_n85_, new_n818_, new_n230_, new_n6081_, new_n317_, new_n746_, new_n399_, new_n2049_, new_n79_, new_n284_, new_n410_, new_n998_, new_n1352_, new_n170_, new_n1007_, new_n669_, new_n2158_, new_n467_, new_n5195_, new_n616_, new_n1559_, new_n205_, new_n1351_, new_n287_, new_n5417_, new_n225_, new_n1501_, y[0], new_n95_, new_n520_, new_n207_, new_n1036_, new_n387_, new_n494_, new_n97_, new_n576_, new_n966_, new_n220_, new_n5687_, new_n648_, new_n5688_, new_n864_, new_n1390_, new_n262_, new_n5850_, new_n471_, new_n522_, new_n367_, new_n486_, new_n541_, new_n678_, new_n148_, new_n649_, new_n405_, new_n2774_, new_n221_, new_n6194_, new_n229_, new_n668_, new_n6291_, new_n161_, new_n1690_, new_n328_, new_n4921_, x[1], new_n5747_, new_n6185_, new_n2859_, new_n448_, new_n2219_, new_n342_, new_n1009_, new_n266_, new_n3287_, new_n231_, new_n419_, new_n246_, new_n3516_, new_n355_, new_n5702_, new_n289_, new_n1168_, new_n1076_, new_n2105_, new_n414_, new_n1536_, new_n350_, new_n1041_, new_n184_, new_n3408_, new_n129_, new_n5058_, new_n715_, new_n751_, new_n149_, new_n1769_, new_n4636_, new_n155_, new_n5713_, new_n370_, new_n2557_, new_n318_, new_n1117_, new_n192_, new_n1309_, new_n354_, new_n1951_, new_n425_, new_n5178_, new_n189_, new_n1603_, new_n159_, new_n617_, new_n1791_, new_n213_, new_n4733_, new_n91_, new_n5786_, new_n6294_, new_n786_, new_n3026_, new_n4973_, new_n979_, new_n1132_, new_n209_, new_n1470_, new_n1222_, new_n3004_, new_n244_, new_n4612_, x[2], new_n339_, new_n509_, new_n495_, new_n4401_, new_n1103_, new_n1641_, new_n481_, new_n2755_, new_n275_, new_n907_, new_n241_, new_n2136_, new_n371_, new_n1922_, new_n169_, new_n611_, new_n271_, new_n1175_, new_n150_, new_n5512_, new_n975_, new_n3025_, new_n214_, new_n5526_, new_n82_, new_n88_, new_n335_, new_n6248_, new_n127_, new_n3122_, new_n460_, new_n3931_, new_n81_, new_n4546_, new_n4632_, new_n378_, new_n3990_, new_n1034_, new_n3541_, new_n243_, new_n5772_, new_n343_, new_n4952_, new_n493_, new_n2188_, new_n153_, new_n735_, new_n164_, new_n5717_, new_n270_, new_n5614_, new_n238_, new_n6074_, new_n383_, new_n1652_, new_n5446_, new_n385_, new_n1243_, new_n269_, new_n869_, new_n179_, new_n5279_, new_n445_, new_n1465_, new_n313_, new_n4570_, new_n465_, new_n5766_, new_n968_, new_n2159_, new_n250_, new_n1463_, new_n204_, new_n5291_, new_n200_, new_n4873_, new_n254_, new_n6202_, new_n676_, new_n4730_, new_n218_, new_n4167_, new_n232_, new_n3575_, new_n2885_, new_n623_, new_n4838_, new_n272_, new_n1514_, new_n701_, new_n3705_, new_n123_, new_n2663_, new_n612_, new_n1133_, new_n224_, new_n5953_, new_n334_, new_n686_, new_n173_, new_n1361_, new_n237_, new_n3218_, new_n183_, new_n2116_, new_n603_, new_n637_, new_n359_, new_n5909_, new_n812_, new_n1137_, new_n2189_, new_n636_, new_n679_, new_n182_, new_n6115_, new_n323_, new_n5795_, new_n151_, new_n1469_, new_n312_, new_n5274_, new_n325_, new_n392_, new_n364_, new_n5311_, new_n324_, new_n5167_})
326'b111??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????110???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????101????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????110?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????? : coef[12] = 1'b0;
326'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[12] = 1'b0;
326'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[12] = 1'b0;
326'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00?? : coef[12] = 1'b0;
326'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[12] = 1'b0;
default : coef[12] = 1'b1;
endcase
casez ({new_n122_, new_n5102_, new_n1093_, new_n2576_, new_n242_, new_n5665_, new_n169_, new_n1739_, new_n225_, new_n5494_, new_n416_, new_n4399_, new_n360_, new_n4168_, new_n220_, new_n5305_, new_n267_, new_n4319_, new_n645_, new_n2504_, new_n463_, new_n3135_, new_n887_, new_n622_, new_n1960_, new_n405_, new_n793_, new_n97_, new_n350_, new_n764_, new_n429_, new_n3378_, new_n219_, new_n1036_, new_n207_, new_n908_, new_n248_, new_n1611_, new_n214_, new_n865_, new_n299_, new_n1602_, new_n356_, new_n5239_, new_n229_, new_n1391_, new_n578_, new_n3266_, new_n6221_, new_n481_, new_n5716_, new_n212_, new_n4380_, new_n378_, new_n3522_, new_n127_, new_n4988_, new_n330_, new_n1385_, new_n897_, new_n1205_, new_n353_, new_n1634_, new_n389_, new_n1645_, new_n469_, new_n5860_, new_n198_, new_n2787_, new_n1792_, new_n121_, new_n5255_, new_n228_, new_n5260_, new_n94_, new_n569_, new_n918_, new_n616_, new_n1065_, new_n488_, new_n2826_, new_n274_, new_n3656_, new_n216_, new_n937_, new_n371_, new_n494_, new_n335_, new_n1228_, new_n524_, new_n2738_, new_n187_, new_n548_, new_n339_, new_n620_, new_n495_, new_n965_, new_n447_, new_n5819_, new_n377_, new_n4355_, new_n1004_, new_n1267_, new_n386_, new_n1727_, new_n530_, new_n1461_, new_n306_, new_n718_, new_n164_, new_n5253_, new_n2368_, new_n179_, new_n5789_, new_n915_, new_n2946_, new_n1825_, new_n2968_, new_n257_, new_n724_, new_n574_, new_n1724_, new_n2877_, new_n2298_, new_n860_, new_n1264_, new_n286_, new_n695_, new_n171_, new_n6019_, new_n564_, new_n643_, new_n6256_, new_n236_, new_n732_, new_n1858_, new_n3132_, new_n168_, new_n2254_, new_n6281_, new_n210_, new_n5399_, new_n2908_, new_n159_, new_n647_, new_n445_, new_n4583_, new_n5962_, new_n6216_, new_n269_, new_n4256_, new_n140_, new_n2661_, new_n279_, new_n1225_, new_n113_, new_n4750_, new_n208_, new_n593_, new_n565_, new_n1363_, new_n1362_, new_n1702_, new_n554_, new_n563_, new_n368_, new_n2067_, new_n310_, new_n990_, new_n151_, new_n1333_, new_n375_, new_n1133_, new_n254_, new_n3225_, new_n132_, new_n5694_, new_n305_, new_n811_, new_n303_, new_n2090_, new_n674_, new_n3699_, new_n312_, new_n3815_, new_n155_, new_n5307_, new_n6289_, new_n1246_, v[2], new_n176_, new_n750_, new_n96_, new_n103_, new_n1122_, new_n213_, new_n2672_, new_n924_, new_n2713_, new_n153_, new_n4896_, new_n517_, new_n982_, new_n158_, new_n4829_, new_n150_, new_n1485_, new_n408_, new_n3589_, new_n265_, new_n5522_, new_n1378_, new_n2521_, new_n202_, new_n3846_, new_n126_, new_n188_, new_n669_, new_n3504_, new_n541_, new_n2659_, new_n170_, new_n5758_, new_n115_, new_n5498_, new_n1177_, new_n1932_, new_n205_, new_n3876_, new_n129_, new_n4362_, new_n253_, new_n675_, new_n401_, new_n854_, new_n157_, new_n5389_, new_n259_, new_n5718_, new_n318_, new_n5010_, new_n765_, new_n2737_, new_n161_, new_n6203_, new_n173_, new_n3144_, new_n123_, new_n1368_, new_n280_, new_n1640_, new_n255_, new_n2282_, new_n546_, new_n1801_, new_n917_, new_n927_, new_n144_, new_n5036_, new_n532_, new_n911_, new_n598_, new_n1152_, new_n145_, new_n5406_, new_n245_, new_n556_, y[2], new_n4611_, new_n542_, new_n2716_, new_n149_, new_n4405_, new_n222_, new_n6095_, new_n243_, new_n1476_, new_n426_, new_n457_, new_n184_, new_n5708_, new_n500_, new_n1901_, new_n438_, new_n657_, new_n272_, new_n4493_, new_n1235_, new_n1986_, new_n300_, new_n2568_, new_n528_, new_n1124_, new_n323_, new_n325_, new_n545_, new_n2520_, new_n722_, new_n2635_, new_n697_, new_n997_, new_n2387_, new_n246_, new_n5382_, new_n162_, new_n5901_, new_n182_, new_n5297_, new_n240_, new_n3722_, new_n716_, new_n1940_, new_n301_, new_n516_, new_n175_, new_n4642_, new_n249_, new_n3405_, new_n275_, new_n1474_, new_n190_, new_n4292_, new_n557_, new_n1023_, new_n293_, new_n3494_, new_n582_, new_n4872_})
328'b10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[13] = 1'b1;
328'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[13] = 1'b1;
328'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[13] = 1'b1;
328'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[13] = 1'b1;
328'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[13] = 1'b1;
default : coef[13] = 1'b0;
endcase
casez ({new_n228_, new_n1595_, new_n142_, new_n1149_, new_n941_, new_n4012_, new_n286_, new_n5339_, new_n299_, new_n1863_, new_n275_, new_n3540_, new_n225_, new_n5880_, new_n171_, new_n4501_, new_n86_, new_n6000_, new_n6128_, new_n281_, new_n521_, new_n164_, new_n3418_, new_n230_, new_n535_, new_n6232_, new_n158_, new_n5756_, new_n1628_, new_n3112_, new_n226_, new_n6066_, new_n552_, new_n3594_, new_n172_, new_n5272_, new_n113_, new_n139_, new_n418_, new_n712_, new_n1059_, new_n170_, new_n1522_, new_n265_, new_n810_, new_n620_, new_n2102_, new_n420_, new_n2738_, new_n116_, new_n232_, new_n126_, new_n409_, new_n511_, new_n1227_, new_n1031_, new_n4281_, new_n551_, new_n5794_, new_n333_, new_n4437_, new_n166_, new_n4127_, new_n5443_, new_n255_, new_n1147_, new_n326_, new_n1454_, new_n312_, new_n752_, new_n223_, new_n6101_, new_n236_, new_n1430_, new_n123_, new_n1342_, new_n1098_, new_n5648_, new_n177_, new_n1140_, new_n217_, new_n1870_, new_n422_, new_n1877_, new_n517_, new_n2158_, new_n648_, new_n2689_, new_n221_, new_n4688_, new_n169_, new_n4981_, new_n340_, new_n3381_, new_n319_, new_n2144_, new_n220_, new_n463_, new_n95_, new_n6078_, new_n387_, new_n4412_, new_n244_, new_n1152_, new_n542_, new_n4226_, new_n403_, new_n442_, new_n214_, new_n5031_, new_n372_, new_n1935_, new_n2311_, new_n388_, new_n3561_, new_n412_, new_n2676_, new_n101_, new_n5859_, new_n229_, new_n2778_, new_n583_, new_n1338_, new_n2903_, new_n1242_, new_n3222_, new_n1788_, new_n484_, new_n4038_, new_n6257_, new_n530_, new_n2702_, new_n279_, new_n3319_, new_n342_, new_n1012_, new_n5447_, new_n159_, new_n4674_, new_n471_, new_n1100_, new_n191_, new_n1457_, new_n215_, new_n1562_, new_n218_, new_n5896_, new_n266_, new_n6204_, v[1], new_n87_, new_n1058_, new_n184_, new_n854_, new_n426_, new_n1071_, new_n175_, new_n977_, new_n1486_, new_n1504_, new_n157_, new_n1533_, new_n174_, new_n4842_, new_n302_, new_n516_, new_n370_, new_n4333_, new_n6162_, new_n283_, new_n960_, new_n2872_, new_n205_, new_n6001_, new_n129_, new_n5257_, new_n396_, new_n612_, new_n185_, new_n4388_, new_n213_, new_n5141_, new_n2108_, new_n4813_, new_n331_, new_n955_, new_n186_, new_n562_, new_n245_, new_n4839_, new_n504_, new_n2047_, new_n350_, new_n812_, new_n515_, new_n673_, new_n1958_, new_n3832_, new_n1547_, new_n2744_, new_n194_, new_n2563_, new_n224_, new_n5461_, new_n267_, new_n4931_, new_n309_, new_n1861_, new_n764_, new_n3500_, new_n481_, new_n1179_, new_n371_, new_n4976_, new_n1494_, new_n2496_, new_n1001_, new_n3564_, new_n100_, new_n768_, new_n781_, new_n310_, new_n1404_, u[1], new_n378_, new_n432_, new_n308_, new_n1835_, new_n250_, new_n1062_, new_n274_, new_n1207_, new_n118_, new_n1045_, new_n451_, new_n4685_, new_n405_, new_n2773_, new_n537_, new_n2700_, x[2], new_n3781_, new_n5924_, new_n677_, new_n1821_, new_n505_, new_n3520_, new_n332_, new_n1211_, new_n287_, new_n986_, new_n122_, new_n5736_, new_n398_, new_n3498_, new_n343_, new_n975_, new_n115_, new_n5809_, new_n381_, new_n2747_, new_n153_, new_n5888_, new_n257_, new_n1201_, new_n94_, new_n130_, new_n769_, new_n386_, new_n1302_, new_n179_, new_n5488_, new_n167_, new_n2293_, new_n151_, new_n4689_, new_n2409_, new_n311_, new_n875_, new_n89_, new_n2828_, new_n375_, new_n424_, new_n269_, new_n5595_, new_n391_, new_n538_, new_n134_, new_n2132_, new_n183_, new_n1051_, new_n293_, new_n4883_, new_n196_, new_n1355_, new_n168_, new_n5838_, new_n647_, new_n3303_, new_n462_, new_n5402_, new_n83_, new_n4992_, new_n182_, new_n6120_, new_n231_, new_n3402_, new_n199_, new_n658_, new_n300_, new_n6027_, new_n144_, new_n4777_, new_n239_, new_n5842_, new_n705_, new_n3272_, new_n148_, new_n222_, new_n993_, new_n6269_, new_n253_, new_n4532_, new_n392_, new_n1757_, new_n2491_, new_n91_, new_n1751_, new_n301_, new_n3956_, new_n98_, new_n3795_, new_n145_, new_n1764_, new_n289_, new_n3634_, new_n318_, new_n5478_, new_n753_, new_n4423_, new_n336_, new_n4895_, new_n258_, new_n1054_, new_n6283_})
345'b11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????110?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110????????????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[14] = 1'b1;
345'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[14] = 1'b1;
345'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??? : coef[14] = 1'b1;
345'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11? : coef[14] = 1'b1;
345'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0 : coef[14] = 1'b1;
default : coef[14] = 1'b0;
endcase
casez ({new_n127_, new_n2095_, new_n286_, new_n821_, new_n6274_, new_n635_, new_n1170_, new_n265_, new_n1075_, new_n2157_, new_n4200_, new_n261_, new_n2607_, new_n179_, new_n5560_, new_n306_, new_n5044_, new_n168_, new_n1026_, new_n373_, new_n4572_, new_n313_, new_n948_, new_n390_, new_n3805_, new_n170_, new_n5542_, new_n6033_, new_n337_, new_n1877_, new_n2503_, new_n4024_, new_n285_, new_n779_, v[0], new_n1445_, new_n305_, new_n4790_, new_n175_, new_n1484_, new_n452_, new_n1041_, new_n713_, new_n3700_, new_n467_, new_n5845_, new_n246_, new_n5620_, new_n409_, new_n525_, new_n166_, new_n4675_, new_n433_, new_n4547_, new_n413_, new_n5762_, new_n157_, new_n1212_, new_n242_, new_n3018_, new_n160_, new_n696_, new_n186_, new_n1278_, new_n85_, new_n5992_, new_n253_, new_n4700_, new_n92_, new_n223_, new_n1680_, new_n241_, new_n2657_, new_n263_, new_n5802_, new_n90_, new_n1206_, new_n1166_, new_n1393_, new_n222_, new_n2671_, new_n397_, new_n961_, new_n178_, new_n5152_, new_n366_, new_n1926_, new_n887_, new_n319_, new_n758_, new_n225_, new_n6114_, new_n277_, new_n5603_, new_n122_, new_n5644_, new_n80_, new_n2798_, new_n382_, new_n1805_, new_n2907_, new_n215_, new_n1768_, new_n583_, new_n4165_, new_n220_, new_n5760_, new_n154_, new_n3013_, new_n486_, new_n1422_, new_n2632_, new_n3560_, new_n340_, new_n4482_, v[2], new_n3311_, new_n162_, new_n5232_, new_n343_, new_n1770_, new_n6150_, new_n2860_, new_n297_, new_n1224_, new_n161_, new_n4761_, new_n2374_, new_n192_, new_n761_, new_n172_, new_n5136_, new_n113_, new_n5473_, new_n1241_, new_n279_, new_n384_, new_n6211_, new_n184_, new_n5634_, new_n218_, new_n591_, new_n332_, new_n1721_, new_n375_, new_n556_, new_n325_, new_n2014_, new_n291_, new_n448_, new_n155_, new_n1139_, new_n355_, new_n675_, new_n478_, new_n2698_, new_n289_, new_n714_, new_n502_, new_n1638_, new_n189_, new_n1915_, new_n190_, new_n4879_, new_n280_, new_n3580_, new_n159_, new_n1007_, new_n256_, new_n1733_, new_n396_, new_n6092_, new_n947_, new_n1547_, new_n210_, new_n773_, new_n145_, new_n5781_, new_n144_, new_n5552_, new_n217_, new_n1462_, new_n1238_, new_n173_, new_n5112_, new_n213_, new_n5903_, new_n185_, new_n672_, new_n255_, new_n1901_, new_n411_, new_n2804_, new_n354_, new_n572_, new_n2437_, new_n350_, new_n717_, new_n407_, new_n1073_, new_n353_, new_n4446_, new_n290_, new_n3283_, new_n1222_, new_n2496_, new_n309_, new_n5052_, new_n163_, new_n3412_, new_n605_, new_n868_, new_n282_, new_n505_, new_n327_, new_n1997_, new_n6237_, new_n198_, new_n4868_, new_n6265_, new_n2867_, new_n4623_, new_n153_, new_n723_, new_n339_, new_n622_, new_n118_, new_n1730_, new_n2098_, new_n606_, new_n3693_, new_n216_, new_n2796_, new_n744_, new_n1942_, new_n142_, new_n5755_, new_n806_, new_n1955_, new_n6254_, new_n211_, new_n4588_, u[0], new_n247_, new_n451_, new_n371_, new_n5206_, new_n1001_, new_n1939_, new_n404_, new_n1581_, new_n495_, new_n620_, new_n121_, new_n1824_, new_n449_, new_n5095_, new_n81_, new_n2681_, new_n389_, new_n1180_, new_n381_, new_n1156_, new_n537_, new_n5325_, new_n317_, new_n711_, new_n1088_, new_n2955_, new_n323_, new_n5811_, new_n171_, new_n6205_, new_n89_, new_n468_, new_n530_, new_n4512_, new_n346_, new_n1037_, new_n151_, new_n4950_, new_n2187_, new_n503_, new_n2161_, new_n266_, new_n859_, new_n1303_, new_n2701_, new_n182_, new_n1457_, new_n344_, new_n866_, new_n251_, new_n1330_, new_n132_, new_n4795_, new_n134_, new_n4523_, new_n238_, new_n563_, new_n199_, new_n5336_, new_n300_, new_n876_, new_n208_, new_n6123_, new_n312_, new_n5097_, new_n200_, new_n2806_, new_n188_, new_n424_, new_n458_, new_n3771_, new_n936_, new_n2819_, new_n782_, new_n1091_, new_n722_, new_n1566_, new_n201_, new_n4366_, new_n167_, new_n1217_, new_n550_, new_n812_, new_n148_, new_n1849_, new_n224_, new_n1055_, new_n123_, new_n3662_, new_n129_, new_n4153_, new_n254_, new_n4016_, new_n293_, new_n2655_, new_n582_, new_n753_, new_n272_, new_n4534_})
342'b10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????00?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[15] = 1'b1;
342'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[15] = 1'b1;
342'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[15] = 1'b1;
default : coef[15] = 1'b0;
endcase
casez ({new_n131_, new_n2989_, new_n765_, new_n5816_, new_n262_, new_n2062_, x[2], new_n264_, new_n387_, new_n377_, new_n863_, new_n2482_, new_n287_, new_n4046_, new_n166_, new_n219_, new_n492_, new_n360_, new_n2722_, new_n169_, new_n1149_, new_n1929_, new_n3614_, new_n648_, new_n1946_, v[2], new_n3991_, new_n520_, new_n522_, new_n221_, new_n5535_, new_n228_, new_n2663_, new_n320_, new_n1908_, new_n225_, new_n1155_, new_n358_, new_n904_, new_n241_, new_n813_, new_n207_, new_n725_, new_n212_, new_n1062_, new_n150_, new_n2717_, new_n388_, new_n1377_, new_n121_, new_n3181_, new_n162_, new_n5210_, new_n211_, new_n5065_, new_n488_, new_n1483_, new_n309_, new_n4780_, new_n115_, new_n3728_, new_n243_, new_n611_, new_n2855_, new_n178_, new_n553_, new_n122_, new_n882_, new_n437_, new_n1434_, new_n328_, new_n865_, new_n83_, new_n220_, new_n412_, new_n6150_, new_n423_, new_n1338_, new_n244_, new_n1839_, new_n5444_, new_n98_, new_n1729_, new_n127_, new_n5313_, new_n1726_, new_n3039_, new_n541_, new_n2827_, new_n154_, new_n1728_, new_n619_, new_n1207_, new_n398_, new_n867_, new_n249_, new_n5905_, new_n509_, new_n601_, new_n330_, new_n3558_, new_n1717_, new_n3315_, new_n1196_, new_n757_, new_n2923_, new_n281_, new_n760_, new_n926_, new_n3341_, new_n311_, new_n2506_, new_n576_, new_n1174_, new_n391_, new_n1186_, new_n137_, new_n6075_, new_n2078_, new_n414_, new_n1535_, new_n192_, new_n468_, new_n1366_, new_n4111_, new_n153_, new_n3473_, new_n439_, new_n4170_, new_n1002_, new_n2519_, new_n88_, new_n580_, new_n6286_, new_n2456_, new_n84_, new_n5214_, new_n197_, new_n2688_, new_n1229_, new_n2697_, new_n307_, new_n5474_, new_n6291_, new_n4661_, new_n97_, new_n920_, new_n1256_, new_n266_, new_n5344_, new_n618_, new_n1039_, new_n167_, new_n231_, new_n728_, new_n218_, new_n1630_, new_n140_, new_n798_, new_n164_, new_n1048_, new_n653_, new_n1884_, new_n2483_, new_n100_, new_n1445_, new_n113_, new_n1218_, new_n172_, new_n4946_, new_n5441_, u[2], new_n4984_, new_n93_, new_n1463_, new_n1577_, new_n1619_, new_n238_, new_n2838_, new_n342_, new_n5954_, v[1], new_n1204_, new_n305_, new_n5388_, new_n194_, new_n3365_, new_n145_, new_n5248_, new_n1793_, new_n181_, new_n3710_, new_n552_, new_n686_, new_n202_, new_n5759_, new_n1750_, new_n4048_, new_n217_, new_n5661_, new_n682_, new_n1880_, new_n438_, new_n1530_, new_n315_, new_n3339_, new_n161_, new_n3444_, new_n213_, new_n5491_, new_n91_, new_n6021_, new_n300_, new_n1469_, new_n129_, new_n858_, new_n334_, new_n1031_, new_n2491_, new_n1205_, new_n5701_, new_n325_, new_n4040_, new_n545_, new_n2635_, new_n6280_, new_n4582_, new_n189_, new_n1359_, new_n422_, new_n688_, new_n259_, new_n1020_, new_n677_, new_n3317_, new_n2387_, new_n296_, new_n2000_, new_n333_, new_n1497_, new_n630_, new_n1341_, new_n157_, new_n1345_, new_n230_, new_n1719_, new_n160_, new_n985_, new_n177_, new_n1323_, new_n185_, new_n3202_, new_n155_, new_n3377_, new_n2063_, new_n2501_, new_n3407_, new_n263_, new_n1840_, new_n5456_, new_n86_, new_n5640_, new_n1247_, new_n335_, new_n4556_, new_n144_, new_n958_, new_n126_, new_n425_, new_n390_, new_n1386_, new_n1710_, new_n3579_, new_n158_, new_n175_, new_n363_, new_n273_, new_n1210_, new_n223_, new_n3304_, new_n2249_, new_n265_, new_n701_, new_n2895_, new_n268_, new_n5124_, new_n500_, new_n1606_, new_n190_, new_n4522_, new_n255_, new_n4922_, new_n515_, new_n1166_, new_n6290_, new_n1019_, new_n2765_, u[0], new_n246_, new_n583_, new_n4581_, new_n326_, new_n995_})
303'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????011?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????110?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??????????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????? : coef[16] = 1'b0;
303'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????? : coef[16] = 1'b0;
303'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??? : coef[16] = 1'b0;
303'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? : coef[16] = 1'b0;
303'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[16] = 1'b0;
default : coef[16] = 1'b1;
endcase
casez ({new_n225_, new_n2591_, new_n267_, new_n5578_, new_n928_, new_n3658_, new_n437_, new_n4279_, new_n755_, new_n3074_, new_n486_, new_n4604_, new_n930_, new_n3599_, new_n604_, new_n2656_, new_n624_, new_n1093_, new_n552_, new_n703_, new_n140_, new_n5545_, new_n166_, new_n573_, new_n160_, new_n1243_, new_n242_, new_n761_, new_n6271_, new_n137_, new_n5324_, new_n580_, new_n1264_, new_n5442_, new_n164_, new_n5890_, new_n286_, new_n1525_, new_n311_, new_n3641_, new_n285_, new_n613_, new_n607_, new_n2159_, new_n178_, new_n1786_, new_n281_, new_n2753_, new_n188_, new_n584_, new_n123_, new_n5304_, new_n305_, new_n1555_, new_n85_, new_n4360_, new_n104_, new_n880_, new_n333_, new_n1142_, new_n296_, new_n4201_, new_n478_, new_n4545_, new_n129_, new_n5946_, new_n325_, new_n1679_, new_n189_, new_n4670_, new_n144_, new_n5817_, new_n186_, new_n2626_, new_n557_, new_n1546_, new_n6239_, new_n153_, new_n352_, new_n1540_, new_n2737_, new_n86_, new_n2823_, new_n502_, new_n4406_, new_n223_, new_n4105_, new_n162_, new_n746_, new_n236_, new_n4701_, new_n641_, new_n1644_, new_n145_, new_n5168_, new_n265_, new_n4676_, new_n170_, new_n1924_, new_n154_, new_n5075_, new_n623_, new_n2707_, new_n387_, new_n1641_, new_n634_, new_n1963_, new_n121_, new_n2395_, new_n553_, new_n3263_, new_n341_, new_n614_, new_n1744_, new_n2522_, new_n194_, new_n5125_, new_n320_, new_n2837_, new_n1005_, new_n2975_, new_n496_, new_n1799_, new_n430_, new_n631_, new_n874_, new_n2940_, new_n227_, new_n4653_, new_n142_, new_n976_, new_n82_, new_n1421_, new_n530_, new_n1022_, new_n2279_, new_n159_, new_n5960_, new_n5922_, new_n210_, new_n1242_, new_n313_, new_n2638_, new_n4595_, new_n132_, new_n463_, new_n179_, new_n5965_, new_n643_, new_n1810_, new_n5925_, new_n350_, new_n368_, new_n485_, new_n3782_, new_n175_, new_n402_, new_n246_, new_n687_, new_n280_, new_n297_, new_n532_, new_n2064_, new_n482_, new_n3173_, new_n256_, new_n534_, new_n84_, new_n3908_, new_n315_, new_n1369_, new_n192_, new_n1356_, new_n272_, new_n5635_, new_n222_, new_n5055_, new_n292_, new_n3666_, new_n239_, new_n911_, new_n90_, new_n954_, new_n318_, new_n1008_, new_n544_, new_n927_, new_n698_, new_n1539_, new_n916_, new_n2963_, new_n277_, new_n5723_, new_n394_, new_n3533_, new_n276_, new_n434_, new_n268_, new_n1449_, new_n263_, new_n2363_, new_n339_, new_n3932_, new_n200_, new_n4018_, new_n271_, new_n4034_, new_n2099_, new_n524_, new_n742_, new_n389_, new_n1635_, new_n81_, new_n3400_, new_n151_, new_n3016_, new_n492_, new_n2595_, new_n615_, new_n1590_, new_n299_, new_n2577_, new_n228_, new_n1980_, new_n244_, new_n1585_, new_n260_, new_n723_, new_n119_, new_n1494_, new_n6265_, new_n1061_, new_n1643_, new_n460_, new_n3776_, new_n904_, new_n923_, new_n508_, new_n1377_, new_n469_, new_n975_, new_n316_, new_n1219_, new_n505_, new_n2942_, new_n405_, new_n3091_, new_n95_, new_n1288_, new_n1063_, new_n3159_, new_n537_, new_n5071_, new_n541_, new_n1157_, new_n356_, new_n980_, new_n473_, new_n5383_, u[0], new_n3683_, new_n447_, new_n1557_, new_n249_, new_n856_, new_n435_, new_n1099_, new_n488_, new_n1732_, new_n330_, new_n4476_, new_n274_, new_n3397_, new_n605_, new_n1610_, new_n711_, new_n3223_, new_n1489_, new_n1804_, new_n381_, new_n4443_, new_n323_, new_n652_, new_n89_, new_n6080_, new_n201_, new_n4104_, new_n88_, new_n5867_, new_n491_, new_n834_, new_n167_, new_n710_, new_n171_, new_n5970_, new_n456_, new_n869_, new_n728_, new_n2706_, new_n218_, new_n827_, new_n214_, new_n4143_, new_n269_, new_n4215_, new_n251_, new_n391_, new_n344_, new_n978_, new_n258_, new_n1582_, new_n373_, new_n5051_, new_n794_, new_n4184_, new_n279_, new_n1745_, new_n1069_, new_n3001_, new_n199_, new_n570_, new_n245_, new_n454_, new_n202_, new_n5165_, new_n303_, new_n627_, new_n208_, new_n849_, new_n334_, new_n355_, new_n433_, new_n4159_, new_n253_, new_n5424_, new_n603_, new_n1625_, new_n1387_, new_n2068_, new_n598_, new_n4782_, new_n1137_, new_n1950_, new_n782_, new_n1548_, new_n157_, new_n4956_, new_n183_, new_n5092_, new_n240_, new_n5968_, new_n1194_, new_n1648_, new_n182_, new_n4678_, new_n411_, new_n4718_, new_n155_, new_n5737_, new_n512_, new_n629_, new_n224_, new_n1516_, new_n1474_, new_n3215_, new_n217_, new_n4004_, new_n531_, new_n2788_, new_n392_, new_n3109_})
371'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[17] = 1'b1;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[17] = 1'b1;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[17] = 1'b1;
default : coef[17] = 1'b0;
endcase
casez ({new_n166_, new_n3635_, new_n122_, new_n1121_, new_n1869_, new_n2913_, new_n480_, new_n5787_, new_n225_, new_n6024_, new_n442_, new_n1177_, new_n368_, new_n4463_, new_n282_, new_n653_, new_n281_, new_n647_, new_n89_, new_n3925_, new_n452_, new_n652_, new_n137_, new_n1589_, new_n261_, new_n1934_, new_n285_, new_n2628_, new_n230_, new_n6122_, new_n164_, new_n5998_, new_n2420_, new_n2904_, new_n134_, new_n4905_, new_n635_, new_n5742_, new_n484_, new_n3364_, new_n342_, new_n1481_, new_n5431_, new_n170_, new_n3847_, new_n6272_, new_n915_, new_n2503_, new_n985_, new_n1267_, new_n552_, new_n1633_, new_n202_, new_n4293_, new_n791_, new_n1661_, new_n278_, new_n854_, new_n232_, new_n964_, new_n103_, new_n661_, u[2], new_n4738_, new_n209_, new_n1890_, new_n321_, new_n2666_, new_n527_, new_n3233_, new_n176_, new_n1410_, new_n434_, new_n497_, new_n672_, new_n3719_, new_n123_, new_n5370_, new_n160_, new_n1146_, new_n242_, new_n596_, new_n340_, new_n3690_, new_n86_, new_n1742_, new_n126_, new_n245_, new_n423_, new_n4889_, new_n169_, new_n3911_, new_n286_, new_n792_, new_n6187_, new_n158_, new_n5242_, new_n467_, new_n3434_, new_n1386_, new_n1884_, new_n264_, new_n2659_, new_n175_, new_n3987_, new_n274_, new_n1559_, new_n517_, new_n5240_, new_n397_, new_n3168_, new_n318_, new_n4997_, new_n221_, new_n1371_, new_n742_, new_n3800_, new_n748_, new_n1635_, new_n561_, new_n1802_, new_n419_, new_n1812_, new_n220_, new_n5615_, new_n788_, new_n999_, new_n384_, new_n2960_, new_n634_, new_n1956_, new_n95_, new_n99_, new_n4667_, new_n244_, new_n5465_, new_n6210_, new_n6284_, new_n437_, new_n2642_, new_n97_, new_n149_, new_n2552_, new_n649_, new_n3049_, new_n553_, new_n3177_, new_n118_, new_n5732_, new_n215_, new_n5073_, new_n247_, new_n5881_, new_n275_, new_n4941_, new_n387_, new_n952_, new_n94_, new_n162_, new_n555_, new_n115_, new_n3869_, new_n4594_, new_n154_, new_n4135_, new_n462_, new_n4282_, new_n269_, new_n2017_, new_n396_, new_n2164_, new_n207_, new_n4291_, new_n192_, new_n6098_, new_n218_, new_n946_, new_n210_, new_n4025_, new_n427_, new_n917_, new_n132_, new_n520_, new_n313_, new_n1254_, new_n171_, new_n6015_, new_n475_, new_n1965_, new_n186_, new_n3102_, new_n161_, new_n5886_, new_n159_, new_n5334_, new_n414_, new_n5705_, new_n433_, new_n5616_, new_n188_, new_n970_, new_n217_, new_n1266_, new_n138_, new_n780_, new_n190_, new_n5353_, new_n184_, new_n910_, new_n222_, new_n1354_, new_n148_, new_n2790_, new_n268_, new_n955_, new_n528_, new_n2847_, new_n157_, new_n5533_, new_n411_, new_n3228_, new_n500_, new_n2735_, new_n205_, new_n1456_, new_n942_, new_n1803_, new_n605_, new_n1948_, new_n821_, new_n4799_, new_n744_, new_n3566_, new_n330_, new_n4402_, new_n524_, new_n1645_, new_n957_, new_n1706_, new_n628_, new_n3904_, new_n262_, new_n1587_, new_n252_, new_n3332_, new_n316_, new_n2843_, new_n287_, new_n2142_, new_n119_, new_n757_, new_n6282_, new_n142_, new_n986_, new_n243_, new_n806_, new_n317_, new_n611_, new_n319_, new_n1617_, new_n204_, new_n5127_, new_n455_, new_n481_, new_n429_, new_n1807_, new_n382_, new_n3801_, new_n377_, new_n798_, new_n153_, new_n1207_, new_n786_, new_n1939_, new_n965_, new_n5082_, new_n582_, new_n2154_, new_n460_, new_n3929_, new_n249_, new_n5509_, new_n638_, new_n1382_, new_n435_, new_n4578_, new_n454_, new_n4891_, new_n602_, new_n1525_, new_n270_, new_n3790_, new_n208_, new_n2153_, new_n336_, new_n2838_, new_n1724_, new_n3229_, new_n346_, new_n6099_, new_n179_, new_n5721_, new_n251_, new_n4692_, new_n140_, new_n3391_, new_n2431_, new_n168_, new_n5539_, new_n642_, new_n3155_, new_n358_, new_n2561_, new_n241_, new_n4613_, new_n289_, new_n627_, new_n380_, new_n4244_, new_n259_, new_n334_, new_n200_, new_n5046_, new_n4831_, new_n253_, new_n1137_, new_n88_, new_n5243_, new_n196_, new_n2667_, new_n201_, new_n2612_, new_n539_, new_n3574_, new_n1586_, new_n3317_, new_n151_, new_n5200_, new_n183_, new_n490_, new_n310_, new_n3496_, new_n301_, new_n840_, new_n182_, new_n637_, new_n240_, new_n5106_, new_n173_, new_n1949_, new_n155_, new_n5973_, new_n145_, new_n5990_, new_n144_, new_n5984_, new_n325_, new_n4202_, new_n6129_, new_n875_, new_n3749_, new_n609_, new_n5387_, new_n199_, new_n1316_, new_n6250_})
366'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[18] = 1'b0;
366'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[18] = 1'b0;
366'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??? : coef[18] = 1'b0;
366'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11? : coef[18] = 1'b0;
366'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0 : coef[18] = 1'b0;
default : coef[18] = 1'b1;
endcase
casez ({new_n221_, new_n3050_, new_n244_, new_n3024_, new_n299_, new_n2722_, new_n659_, new_n1929_, new_n487_, new_n1597_, new_n247_, new_n5281_, new_n360_, new_n1921_, new_n6268_, new_n223_, new_n4986_, new_n160_, new_n5096_, new_n220_, new_n726_, new_n416_, new_n3489_, new_n267_, new_n5517_, new_n770_, new_n6127_, new_n435_, new_n3298_, new_n127_, new_n4524_, new_n341_, new_n1351_, new_n767_, new_n2505_, new_n121_, new_n665_, new_n650_, new_n2780_, new_n262_, new_n4089_, new_n492_, new_n5193_, new_n2883_, new_n471_, new_n3668_, new_n216_, new_n4779_, new_n212_, new_n1600_, new_n1179_, new_n4212_, new_n310_, new_n634_, new_n387_, new_n2970_, new_n437_, new_n614_, new_n350_, new_n5677_, new_n194_, new_n4047_, new_n6195_, new_n377_, new_n3040_, new_n6253_, new_n353_, new_n5205_, new_n2245_, new_n6294_, new_n95_, new_n4601_, new_n430_, new_n949_, new_n81_, new_n275_, new_n308_, new_n131_, new_n5803_, new_n142_, new_n1153_, new_n97_, new_n1729_, u[1], new_n207_, new_n481_, new_n786_, new_n3535_, new_n460_, new_n2747_, new_n293_, new_n789_, new_n122_, new_n3734_, new_n1581_, new_n3746_, new_n493_, new_n1207_, new_n271_, new_n4414_, new_n442_, new_n554_, new_n260_, new_n611_, new_n83_, new_n5421_, new_n214_, new_n1211_, new_n82_, new_n1900_, new_n395_, new_n3380_, new_n153_, new_n986_, new_n257_, new_n601_, new_n671_, new_n1049_, new_n537_, new_n1630_, new_n330_, new_n404_, new_n211_, new_n1360_, new_n103_, new_n1582_, new_n104_, new_n4910_, new_n2456_, new_n171_, new_n798_, new_n6130_, new_n305_, new_n1243_, x[2], new_n88_, new_n626_, new_n391_, new_n6065_, new_n166_, new_n5358_, new_n2877_, new_n4584_, new_n158_, new_n978_, new_n926_, new_n1372_, new_n226_, new_n4090_, new_n134_, new_n646_, new_n132_, new_n2304_, new_n446_, new_n1775_, new_n6272_, new_n179_, new_n5693_, new_n2870_, new_n168_, new_n1329_, new_n270_, new_n747_, new_n137_, new_n370_, new_n417_, new_n159_, new_n1860_, new_n427_, new_n5256_, new_n414_, new_n5151_, new_n210_, new_n4631_, new_n285_, new_n1089_, new_n683_, new_n1039_, new_n187_, new_n4924_, new_n224_, new_n6068_, new_n321_, new_n1463_, new_n1230_, new_n208_, new_n5393_, new_n703_, new_n4039_, new_n301_, new_n1106_, new_n313_, new_n5303_, new_n238_, new_n1169_, new_n140_, new_n6088_, new_n218_, new_n5599_, new_n324_, new_n5026_, new_n196_, new_n2339_, new_n199_, new_n311_, y[2], new_n1204_, new_n1477_, new_n246_, new_n963_, new_n157_, new_n1631_, new_n126_, new_n232_, new_n6251_, new_n259_, new_n5709_, new_n282_, new_n982_, new_n557_, new_n2759_, new_n189_, new_n1573_, new_n317_, new_n2666_, new_n240_, new_n1627_, new_n230_, new_n2690_, new_n528_, new_n870_, new_n175_, new_n755_, new_n303_, new_n1113_, new_n855_, new_n1400_, new_n242_, new_n2612_, new_n177_, new_n5637_, new_n145_, new_n1383_, new_n433_, new_n1027_, new_n1214_, new_n2936_, new_n743_, new_n5222_, new_n641_, new_n1016_, new_n213_, new_n5764_, new_n1576_, new_n3099_, new_n170_, new_n2066_, new_n682_, new_n4900_, new_n184_, new_n2124_, new_n149_, new_n4409_, new_n1550_, new_n2571_, new_n426_, new_n5034_, new_n268_, new_n272_, new_n190_, new_n5348_, new_n539_, new_n4214_, new_n161_, new_n6013_, new_n255_, new_n1524_, new_n2909_, new_n1475_, new_n1796_, new_n1166_, new_n1951_, new_n186_, new_n4162_, new_n90_, new_n5009_, new_n222_, new_n520_, new_n515_, new_n984_, new_n422_, new_n3300_, new_n250_, new_n2705_, new_n173_, new_n5489_, new_n2871_, new_n204_, new_n1217_, new_n144_, new_n5192_, new_n490_, new_n1133_, x[1], new_n2112_, new_n155_, new_n5561_, new_n708_, new_n1394_, new_n217_, new_n858_, new_n1803_, new_n4527_, new_n478_, new_n2623_, new_n89_, new_n1300_, new_n502_, new_n3512_, new_n183_, new_n1708_, new_n245_, new_n5224_, new_n791_, new_n1182_, new_n582_, new_n960_, new_n1137_, new_n1648_, new_n697_, new_n2126_, u[2], new_n182_, new_n202_, new_n679_, new_n2757_, new_n906_, new_n3592_})
338'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????? : coef[19] = 1'b0;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????? : coef[19] = 1'b0;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111???? : coef[19] = 1'b0;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[19] = 1'b0;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[19] = 1'b0;
default : coef[19] = 1'b1;
endcase
casez ({new_n228_, new_n5471_, new_n225_, new_n2113_, new_n493_, new_n1068_, new_n247_, new_n3646_, new_n221_, new_n685_, new_n429_, new_n3539_, new_n161_, new_n816_, new_n131_, new_n5936_, new_n282_, new_n634_, new_n2434_, new_n1544_, new_n5282_, new_n668_, new_n766_, new_n6287_, new_n360_, new_n3388_, new_n1504_, new_n3756_, new_n191_, new_n1753_, new_n341_, new_n1435_, new_n952_, new_n1881_, new_n2461_, new_n215_, new_n1272_, y[0], new_n97_, new_n1005_, new_n295_, new_n1344_, new_n2311_, new_n404_, new_n3357_, new_n248_, new_n3615_, new_n496_, new_n6096_, new_n162_, new_n4713_, new_n126_, new_n2146_, new_n98_, new_n323_, new_n966_, new_n898_, new_n3290_, new_n343_, new_n605_, new_n537_, new_n4035_, new_n327_, new_n3584_, new_n79_, new_n84_, new_n2843_, new_n723_, new_n1804_, new_n121_, new_n4754_, new_n127_, new_n859_, new_n495_, new_n790_, new_n154_, new_n725_, new_n150_, new_n4977_, new_n907_, new_n3316_, new_n139_, new_n5218_, new_n389_, new_n4210_, new_n2098_, new_n216_, new_n5000_, new_n212_, new_n5544_, x[1], new_n2800_, new_n214_, new_n3037_, new_n194_, new_n735_, new_n243_, new_n1471_, new_n1063_, new_n3720_, new_n480_, new_n4031_, new_n118_, new_n5084_, new_n447_, new_n3841_, new_n115_, new_n1431_, new_n353_, new_n3926_, new_n249_, new_n5638_, new_n258_, new_n3859_, new_n430_, new_n1473_, new_n381_, new_n4462_, new_n633_, new_n4176_, new_n505_, new_n3778_, new_n116_, new_n3412_, new_n388_, new_n3396_, new_n524_, new_n583_, new_n164_, new_n5484_, new_n230_, new_n5655_, new_n176_, new_n4940_, new_n140_, new_n3448_, new_n218_, new_n1828_, new_n160_, new_n593_, new_n445_, new_n1870_, new_n313_, new_n1027_, new_n226_, new_n5059_, new_n604_, new_n5229_, new_n930_, new_n2701_, new_n311_, new_n1626_, new_n6044_, new_n624_, new_n3009_, new_n2465_, new_n178_, new_n5470_, new_n137_, new_n4531_, new_n448_, new_n1224_, new_n6220_, new_n6281_, new_n192_, new_n5365_, new_n5454_, new_n134_, new_n5851_, new_n367_, new_n2109_, new_n4640_, new_n386_, new_n2729_, new_n391_, new_n751_, new_n276_, new_n462_, new_n174_, new_n1897_, new_n454_, new_n4901_, new_n270_, new_n4182_, new_n132_, new_n1612_, new_n2085_, new_n538_, new_n912_, new_n88_, new_n1220_, new_n179_, new_n5971_, new_n1464_, new_n2515_, new_n439_, new_n1722_, new_n393_, new_n1468_, new_n151_, new_n2339_, new_n503_, new_n5250_, new_n269_, new_n679_, new_n373_, new_n676_, new_n224_, new_n6138_, new_n535_, new_n2983_, new_n187_, new_n1556_, new_n306_, new_n3329_, new_n241_, new_n2561_, new_n199_, new_n6112_, new_n171_, new_n5914_, new_n281_, new_n510_, x[2], new_n101_, new_n617_, new_n305_, new_n808_, new_n173_, new_n5503_, new_n253_, new_n5666_, new_n312_, new_n4811_, new_n278_, new_n2683_, new_n452_, new_n812_, new_n104_, new_n586_, new_n232_, new_n3874_, new_n155_, new_n5898_, new_n418_, new_n2733_, new_n177_, new_n5538_, new_n413_, new_n5285_, new_n717_, new_n943_, new_n354_, new_n1129_, new_n992_, new_n2128_, new_n545_, new_n3701_, new_n458_, new_n1113_, new_n202_, new_n5678_, new_n145_, new_n423_, new_n236_, new_n3751_, new_n263_, new_n5897_, new_n245_, new_n1893_, new_n1019_, new_n1393_, new_n715_, new_n3998_, new_n109_, new_n2801_, new_n275_, new_n1736_, new_n170_, new_n5932_, new_n175_, new_n5895_, new_n302_, new_n1491_, new_n365_, new_n608_, new_n297_, new_n355_, new_n159_, new_n811_, new_n210_, new_n2691_, new_n1191_, new_n1642_, new_n272_, new_n4719_, new_n217_, new_n5627_, new_n318_, new_n5013_, new_n184_, new_n5680_, new_n333_, new_n1901_, new_n144_, new_n5309_, new_n268_, new_n3973_, new_n222_, new_n1895_, new_n239_, new_n5741_, new_n205_, new_n1754_, new_n289_, new_n5179_, new_n186_, new_n3613_, new_n984_, new_n4396_, new_n673_, new_n4415_, new_n467_, new_n1917_, new_n594_, new_n3069_, new_n981_, new_n1091_, new_n2189_, new_n123_, new_n5531_, new_n450_, new_n1668_, new_n1548_, new_n2813_, new_n409_, new_n3478_, new_n246_, new_n1772_, new_n183_, new_n4343_, new_n153_, new_n6118_, new_n344_, new_n5172_, new_n356_, new_n1849_, new_n190_, new_n5884_, new_n931_, new_n5724_, new_n204_, new_n4149_, new_n189_, new_n5060_, new_n325_, new_n995_, new_n238_, new_n1834_, new_n280_, new_n2103_, new_n89_, new_n3899_, new_n347_, new_n5600_, new_n129_, new_n5287_})
367'b10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????111??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????001????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[20] = 1'b1;
367'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????? : coef[20] = 1'b1;
367'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[20] = 1'b1;
367'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[20] = 1'b1;
367'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[20] = 1'b1;
default : coef[20] = 1'b0;
endcase
casez ({new_n713_, new_n1622_, new_n219_, new_n4083_, new_n262_, new_n2643_, new_n764_, new_n2619_, new_n943_, new_n2632_, new_n309_, new_n2656_, new_n267_, new_n5893_, new_n974_, new_n3239_, new_n220_, new_n4051_, new_n480_, new_n1119_, new_n416_, new_n2689_, new_n1889_, new_n3609_, new_n225_, new_n2395_, new_n283_, new_n442_, new_n6049_, new_n367_, new_n499_, new_n103_, new_n4913_, new_n165_, new_n4229_, new_n244_, new_n5799_, new_n405_, new_n3913_, new_n95_, new_n5710_, new_n345_, new_n1344_, new_n94_, new_n1254_, new_n277_, new_n3537_, new_n331_, new_n4431_, new_n228_, new_n6111_, new_n127_, new_n6193_, new_n268_, new_n5176_, new_n461_, new_n821_, new_n351_, new_n2615_, new_n2625_, new_n2774_, new_n504_, new_n1704_, new_n139_, new_n976_, new_n1671_, new_n4576_, new_n631_, new_n4473_, new_n898_, new_n3200_, new_n366_, new_n460_, new_n122_, new_n1136_, new_n324_, new_n5327_, new_n330_, new_n1651_, new_n776_, new_n1634_, new_n505_, new_n1389_, new_n151_, new_n988_, new_n531_, new_n2563_, new_n360_, new_n4037_, new_n221_, new_n1384_, new_n290_, new_n4492_, new_n169_, new_n1730_, new_n153_, new_n2793_, new_n6230_, new_n308_, new_n3596_, new_n249_, new_n5134_, new_n275_, new_n1723_, new_n82_, new_n99_, new_n3318_, new_n251_, new_n2778_, new_n115_, new_n1483_, new_n1920_, new_n4235_, new_n327_, new_n1398_, new_n250_, new_n1861_, new_n1580_, new_n3871_, new_n353_, new_n4196_, new_n321_, new_n937_, new_n958_, new_n4376_, new_n1579_, new_n4179_, y[1], new_n449_, new_n469_, new_n241_, new_n881_, new_n744_, new_n3521_, new_n389_, new_n2747_, new_n712_, new_n1489_, new_n1935_, new_n4484_, new_n633_, new_n638_, new_n435_, new_n537_, new_n494_, new_n1798_, new_n340_, new_n3862_, new_n162_, new_n711_, new_n142_, new_n5887_, new_n680_, new_n3257_, new_n473_, new_n620_, new_n121_, new_n264_, new_n347_, new_n281_, new_n1242_, new_n311_, new_n551_, new_n171_, new_n5749_, new_n270_, new_n3894_, new_n140_, new_n4808_, new_n176_, new_n4968_, new_n166_, new_n626_, new_n179_, new_n6147_, new_n160_, new_n5752_, new_n1578_, new_n3587_, new_n194_, new_n1349_, new_n375_, new_n5227_, new_n368_, new_n4715_, new_n164_, new_n5277_, new_n158_, new_n6005_, new_n132_, new_n948_, new_n137_, new_n5008_, new_n261_, new_n4315_, new_n266_, new_n5839_, new_n313_, new_n779_, new_n2884_, new_n168_, new_n5844_, new_n682_, new_n1577_, new_n2406_, new_n1002_, new_n1163_, new_n297_, new_n3594_, new_n393_, new_n3475_, new_n210_, new_n3616_, new_n414_, new_n652_, new_n106_, new_n260_, new_n2543_, new_n391_, new_n970_, new_n2906_, new_n3416_, new_n5450_, new_n2842_, new_n2951_, new_n307_, new_n5540_, new_n419_, new_n439_, new_n3419_, new_n279_, new_n1089_, new_n342_, new_n562_, new_n4608_, new_n184_, new_n1243_, new_n2899_, new_n191_, new_n4023_, new_n248_, new_n2605_, new_n89_, new_n819_, new_n535_, new_n656_, new_n2085_, new_n306_, new_n4080_, new_n88_, new_n1876_, new_n113_, new_n5360_, new_n547_, new_n1813_, new_n167_, new_n1749_, new_n703_, new_n1039_, new_n237_, new_n784_, new_n1220_, new_n2931_, new_n187_, new_n577_, new_n441_, new_n1652_, new_n285_, new_n1069_, new_n445_, new_n2140_, new_n305_, new_n617_, new_n273_, new_n2608_, new_n155_, new_n1896_, new_n272_, new_n4061_, new_n284_, new_n482_, new_n129_, new_n1727_, new_n630_, new_n837_, new_n173_, new_n1565_, new_n157_, new_n5875_, new_n177_, new_n5824_, new_n175_, new_n5537_, new_n92_, new_n5587_, new_n86_, new_n1007_, new_n123_, new_n2001_, new_n394_, new_n3570_, new_n85_, new_n6072_, new_n586_, new_n1101_, new_n286_, new_n5566_, new_n500_, new_n644_, new_n930_, new_n1018_, new_n390_, new_n2158_, new_n410_, new_n5234_, new_n2650_, new_n2944_, new_n178_, new_n2555_, new_n148_, new_n3110_, new_n536_, new_n5646_, new_n253_, new_n3845_, new_n354_, new_n747_, new_n256_, new_n5173_, new_n217_, new_n1684_, new_n280_, new_n5216_, new_n2172_, new_n292_, new_n303_, new_n213_, new_n5590_, new_n222_, new_n561_, new_n498_, new_n2611_, new_n189_, new_n4967_, new_n4636_, new_n150_, new_n2114_, new_n246_, new_n5130_, new_n672_, new_n872_, new_n318_, new_n737_, new_n215_, new_n1841_, new_n502_, new_n1167_, new_n190_, new_n1715_, new_n478_, new_n1480_, y[2], new_n87_, new_n1476_, new_n146_, new_n4648_, new_n240_, new_n900_, new_n350_, new_n704_, new_n763_, new_n2813_, new_n144_, new_n3898_, new_n323_, new_n5462_, new_n467_, new_n795_, new_n334_, new_n2399_, new_n612_, new_n2104_, new_n450_, new_n3507_, new_n346_, new_n1718_, new_n325_, new_n2024_, new_n316_, new_n1474_, new_n204_, new_n5117_, new_n202_, new_n1134_, new_n6252_, new_n715_, new_n1619_, new_n205_, new_n1215_, new_n238_, new_n5593_, new_n254_, new_n1428_, new_n312_, new_n3127_})
405'b11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????101?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00?????????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????? : coef[21] = 1'b0;
405'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[21] = 1'b0;
405'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[21] = 1'b0;
405'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[21] = 1'b0;
405'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[21] = 1'b0;
default : coef[21] = 1'b1;
endcase
casez ({new_n179_, new_n5318_, new_n410_, new_n2507_, new_n175_, new_n1558_, new_n157_, new_n5843_, new_n284_, new_n1208_, new_n713_, new_n5707_, new_n278_, new_n1516_, new_n247_, new_n1595_, new_n228_, new_n1026_, new_n164_, new_n3696_, new_n2368_, new_n176_, new_n468_, x[0], new_n261_, new_n1029_, new_n306_, new_n1828_, new_n160_, new_n6199_, new_n280_, new_n4204_, new_n230_, new_n1438_, new_n101_, new_n3637_, new_n189_, new_n5885_, new_n420_, new_n3336_, new_n213_, new_n1118_, new_n158_, new_n1659_, new_n225_, new_n6116_, new_n262_, new_n2157_, new_n619_, new_n2656_, new_n198_, new_n724_, new_n5433_, new_n2465_, new_n218_, new_n5820_, new_n1251_, new_n408_, new_n3530_, new_n265_, new_n484_, new_n375_, new_n4575_, new_n1037_, new_n3129_, new_n427_, new_n624_, new_n236_, new_n5123_, new_n643_, new_n774_, new_n488_, new_n1209_, new_n145_, new_n5573_, new_n178_, new_n3244_, new_n1395_, new_n3823_, new_n124_, new_n3031_, new_n318_, new_n2058_, new_n123_, new_n5571_, new_n967_, new_n1898_, new_n272_, new_n4716_, new_n797_, new_n1082_, new_n239_, new_n1453_, new_n613_, new_n3281_, new_n170_, new_n814_, new_n240_, new_n3169_, new_n246_, new_n4917_, new_n416_, new_n4219_, new_n282_, new_n2654_, new_n220_, new_n1368_, new_n269_, new_n322_, new_n6257_, new_n172_, new_n946_, new_n171_, new_n1669_, new_n747_, new_n1629_, new_n414_, new_n1191_, new_n159_, new_n6069_, new_n302_, new_n702_, new_n161_, new_n617_, new_n370_, new_n4784_, new_n192_, new_n2224_, new_n2883_, new_n4586_, new_n463_, new_n4358_, new_n384_, new_n3034_, new_n766_, new_n1104_, new_n94_, new_n614_, new_n127_, new_n4078_, new_n113_, new_n2299_, new_n4643_, new_n279_, new_n762_, new_n205_, new_n5664_, new_n283_, new_n3975_, new_n185_, new_n5430_, new_n202_, new_n4729_, new_n422_, new_n916_, new_n188_, new_n331_, new_n169_, new_n3645_, new_n874_, new_n4479_, new_n249_, new_n3687_, new_n295_, new_n2583_, new_n207_, new_n631_, new_n442_, new_n3560_, new_n309_, new_n5769_, new_n555_, new_n3712_, new_n650_, new_n807_, new_n299_, new_n4851_, new_n142_, new_n1862_, new_n96_, new_n579_, new_n706_, new_n522_, new_n2745_, new_n229_, new_n1768_, new_n451_, new_n1344_, new_n373_, new_n1902_, new_n556_, new_n877_, new_n106_, new_n1003_, new_n2899_, new_n1624_, new_n3275_, new_n315_, new_n1715_, new_n350_, new_n1625_, new_n500_, new_n2729_, new_n382_, new_n3949_, new_n426_, new_n1430_, new_n184_, new_n3211_, new_n1096_, new_n1603_, new_n91_, new_n657_, new_n90_, new_n95_, new_n1601_, x[2], new_n316_, new_n578_, new_n82_, new_n1361_, new_n290_, new_n3735_, new_n1047_, new_n1159_, new_n139_, new_n2130_, new_n300_, new_n5547_, new_n2442_, new_n776_, new_n4309_, new_n98_, new_n181_, new_n524_, new_n313_, new_n566_, new_n200_, new_n3828_, new_n1850_, new_n2161_, new_n391_, new_n603_, new_n311_, new_n4898_, new_n462_, new_n2000_, new_n445_, new_n1855_, new_n1566_, new_n3259_, new_n140_, new_n3206_, new_n259_, new_n2764_, new_n355_, new_n5359_, new_n399_, new_n1042_, new_n89_, new_n4914_, new_n602_, new_n1449_, new_n263_, new_n692_, new_n334_, new_n4015_, new_n336_, new_n533_, new_n173_, new_n5188_, new_n1545_, new_n2823_, new_n208_, new_n1083_, new_n727_, new_n997_, new_n190_, new_n2749_, new_n324_, new_n2416_, new_n103_, new_n757_, new_n121_, new_n2132_, new_n1781_, new_n2867_, new_n809_, new_n1643_, new_n194_, new_n5730_, new_n509_, new_n980_, new_n417_, new_n1213_, new_n6279_, new_n616_, new_n1725_, new_n154_, new_n4791_, new_n1142_, new_n1382_, new_n250_, new_n2309_, new_n604_, new_n1063_, new_n5439_, new_n541_, new_n1472_, new_n134_, new_n5996_, new_n214_, new_n4497_, new_n368_, new_n679_, new_n5438_, new_n301_, new_n626_, new_n167_, new_n778_, new_n237_, new_n5790_, new_n232_, new_n3203_, new_n129_, new_n5878_, new_n325_, new_n869_, new_n222_, new_n1348_, new_n182_, new_n750_, new_n346_, new_n595_, new_n274_, new_n867_, new_n459_, new_n1404_, new_n639_, new_n1872_, new_n389_, new_n2839_, new_n2367_, new_n131_, new_n693_, new_n216_, new_n4478_, new_n271_, new_n4447_, new_n133_, new_n4848_, new_n341_, new_n1607_, new_n162_, new_n856_, new_n83_, new_n5943_, new_n132_, new_n4008_, new_n224_, new_n1464_, new_n204_, new_n909_, new_n6231_, new_n293_, new_n637_, new_n545_, new_n3458_, new_n186_, new_n4794_, new_n254_, new_n1912_, new_n289_, new_n1110_, new_n187_, new_n705_})
376'b10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????101????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[22] = 1'b1;
376'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[22] = 1'b1;
376'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[22] = 1'b1;
376'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[22] = 1'b1;
376'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[22] = 1'b1;
default : coef[22] = 1'b0;
endcase
casez ({new_n551_, new_n1928_, v[1], new_n299_, new_n871_, new_n176_, new_n2996_, new_n139_, new_n5230_, new_n522_, new_n3487_, new_n221_, new_n4856_, new_n220_, new_n755_, new_n223_, new_n1574_, new_n262_, new_n1206_, new_n416_, new_n635_, new_n247_, new_n5316_, new_n122_, new_n1218_, new_n648_, new_n4140_, new_n244_, new_n4351_, new_n372_, new_n1961_, new_n822_, new_n994_, new_n405_, new_n721_, new_n487_, new_n788_, new_n764_, new_n5384_, y[0], new_n698_, new_n1013_, new_n4223_, new_n81_, new_n5692_, new_n267_, new_n916_, new_n82_, new_n2586_, new_n442_, new_n751_, new_n6032_, new_n541_, new_n1375_, new_n619_, new_n3527_, new_n493_, new_n2588_, u[0], new_n1195_, new_n3347_, new_n6276_, new_n214_, new_n4982_, new_n169_, new_n5941_, new_n320_, new_n2745_, new_n6221_, new_n495_, new_n742_, new_n142_, new_n3839_, new_n447_, new_n1647_, new_n143_, new_n757_, new_n371_, new_n2998_, x[1], new_n3941_, new_n150_, new_n1472_, new_n606_, new_n3843_, new_n271_, new_n5852_, new_n381_, new_n1181_, new_n211_, new_n1471_, new_n356_, new_n2004_, new_n5444_, new_n335_, new_n1035_, new_n249_, new_n867_, new_n293_, new_n5379_, new_n1001_, new_n4390_, new_n339_, new_n2732_, new_n620_, new_n1034_, new_n290_, new_n749_, new_n453_, new_n579_, new_n207_, new_n601_, new_n131_, new_n4348_, new_n241_, new_n1489_, new_n524_, new_n3541_, new_n1249_, new_n605_, new_n2966_, new_n389_, new_n583_, new_n154_, new_n3273_, new_n379_, new_n1224_, new_n270_, new_n855_, new_n278_, new_n6191_, new_n235_, new_n1370_, new_n565_, new_n2969_, new_n137_, new_n4963_, new_n525_, new_n1174_, new_n484_, new_n3477_, new_n166_, new_n521_, new_n134_, new_n1010_, new_n784_, new_n3148_, new_n386_, new_n1933_, new_n168_, new_n1383_, new_n610_, new_n992_, new_n158_, new_n1200_, new_n112_, new_n2645_, new_n113_, new_n5392_, v[0], new_n1444_, new_n2884_, new_n5448_, new_n4594_, new_n159_, new_n6082_, new_n161_, new_n468_, new_n368_, new_n396_, new_n192_, new_n760_, new_n445_, new_n5317_, new_n313_, new_n5997_, new_n138_, new_n2842_, new_n285_, new_n471_, new_n132_, new_n5626_, new_n391_, new_n4218_, new_n191_, new_n547_, new_n269_, new_n4285_, new_n385_, new_n2293_, new_n300_, new_n577_, new_n86_, new_n243_, new_n990_, new_n200_, new_n568_, new_n172_, new_n2633_, new_n6267_, new_n196_, new_n1562_, new_n5437_, new_n88_, new_n5201_, new_n179_, new_n1846_, new_n171_, new_n5972_, new_n311_, new_n1553_, new_n2297_, new_n151_, new_n2869_, new_n810_, new_n1194_, new_n182_, new_n695_, new_n342_, new_n3373_, new_n266_, new_n2622_, new_n204_, new_n4459_, new_n456_, new_n1134_, new_n441_, new_n1343_, new_n306_, new_n4629_, new_n254_, new_n1037_, new_n373_, new_n2179_, new_n186_, new_n3070_, new_n281_, new_n696_, new_n303_, new_n584_, new_n129_, new_n5408_, new_n291_, new_n713_, new_n104_, new_n518_, new_n250_, new_n3481_, new_n1543_, new_n1898_, new_n500_, new_n5466_, new_n230_, new_n5343_, new_n123_, new_n4156_, new_n315_, new_n2711_, new_n458_, new_n1129_, new_n177_, new_n3278_, new_n144_, new_n340_, new_n259_, new_n2521_, new_n6261_, new_n1071_, new_n1885_, new_n3704_, new_n236_, new_n5209_, new_n178_, new_n586_, new_n399_, new_n1397_, new_n289_, new_n4904_, new_n170_, new_n1741_, new_n325_, new_n501_, new_n476_, new_n981_, new_n297_, new_n1486_, new_n302_, new_n2655_, new_n414_, new_n5549_, new_n280_, new_n322_, new_n155_, new_n5611_, new_n205_, new_n767_, new_n1057_, new_n4211_, new_n924_, new_n2118_, new_n715_, new_n4453_, new_n463_, new_n1539_, new_n90_, new_n2334_, new_n217_, new_n1500_, new_n275_, new_n2114_, new_n426_, new_n1053_, new_n268_, new_n1387_, new_n502_, new_n1423_, new_n246_, new_n440_, new_n174_, new_n1748_, new_n328_, new_n1475_, new_n433_, new_n2736_, new_n434_, new_n504_, y[2], new_n420_, new_n602_, new_n334_, new_n3766_, new_n450_, new_n1699_, new_n1038_, new_n1205_, new_n208_, new_n861_, new_n424_, new_n457_, new_n222_, new_n4774_, new_n438_, new_n1225_, new_n336_, new_n1135_, new_n324_, new_n539_, new_n157_, new_n5184_, new_n2126_, new_n2836_, new_n173_, new_n5944_, new_n358_, new_n2705_, new_n167_, new_n2558_, new_n145_, new_n5879_, new_n529_, new_n873_, new_n148_, new_n346_, new_n428_, new_n232_, new_n1040_, new_n263_, new_n1407_, new_n194_, new_n4912_, new_n187_, new_n6017_, new_n365_, new_n2773_, new_n199_, new_n727_, new_n258_, new_n5948_})
378'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????001????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????? : coef[23] = 1'b0;
378'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[23] = 1'b0;
378'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110?????????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[23] = 1'b0;
378'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[23] = 1'b0;
378'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10 : coef[23] = 1'b0;
default : coef[23] = 1'b1;
endcase
casez ({new_n230_, new_n5959_, new_n480_, new_n3170_, new_n405_, new_n497_, new_n942_, new_n1814_, new_n228_, new_n4283_, new_n221_, new_n6100_, new_n265_, new_n5649_, new_n2151_, new_n3297_, new_n2654_, new_n3565_, new_n1385_, new_n1960_, new_n299_, new_n3995_, y[2], new_n135_, new_n1338_, new_n742_, new_n2582_, new_n192_, new_n5323_, new_n1266_, new_n2517_, new_n121_, new_n4539_, new_n283_, new_n2741_, new_n220_, new_n4932_, new_n127_, new_n5645_, new_n95_, new_n5653_, new_n492_, new_n777_, new_n244_, new_n758_, new_n486_, new_n698_, new_n310_, new_n5679_, new_n1170_, new_n4573_, new_n98_, new_n277_, new_n2916_, new_n372_, new_n4486_, new_n262_, new_n5320_, new_n149_, new_n4694_, new_n250_, new_n1376_, new_n207_, new_n4850_, new_n79_, new_n2798_, new_n522_, new_n1735_, new_n435_, new_n632_, new_n864_, new_n952_, new_n215_, new_n4146_, new_n2677_, new_n4989_, new_n194_, new_n4987_, new_n335_, new_n748_, new_n216_, new_n5087_, new_n1202_, new_n3301_, new_n282_, new_n3698_, new_n378_, new_n3714_, new_n2442_, new_n97_, new_n4878_, new_n122_, new_n150_, new_n201_, new_n345_, new_n987_, new_n107_, new_n167_, new_n416_, new_n212_, new_n1150_, new_n341_, new_n2704_, new_n6237_, new_n267_, new_n1021_, new_n162_, new_n5235_, new_n214_, new_n1061_, new_n935_, new_n1623_, new_n169_, new_n4978_, new_n5449_, new_n495_, new_n5226_, new_n616_, new_n907_, new_n249_, new_n5807_, new_n225_, new_n4373_, new_n604_, new_n5138_, new_n1001_, new_n1610_, new_n950_, new_n1404_, new_n1872_, new_n4472_, new_n1706_, new_n2839_, new_n275_, new_n711_, new_n241_, new_n2723_, new_n131_, new_n5128_, new_n6236_, new_n330_, new_n749_, new_n473_, new_n798_, new_n305_, new_n860_, new_n462_, new_n964_, new_n137_, new_n5835_, new_n2494_, new_n446_, new_n552_, new_n218_, new_n718_, new_n164_, new_n2055_, new_n166_, new_n1088_, new_n176_, new_n3524_, new_n373_, new_n3860_, new_n177_, new_n978_, new_n86_, new_n5157_, new_n6130_, new_n142_, new_n4869_, new_n386_, new_n4125_, new_n6031_, new_n445_, new_n4749_, new_n286_, new_n1292_, new_n306_, new_n5499_, new_n139_, new_n1059_, new_n178_, new_n4837_, new_n171_, new_n5633_, new_n368_, new_n448_, new_n1169_, new_n4197_, new_n140_, new_n2267_, new_n2078_, new_n4618_, new_n159_, new_n5299_, new_n5926_, new_n210_, new_n4344_, new_n970_, new_n1174_, new_n342_, new_n946_, new_n113_, new_n3729_, new_n901_, new_n3934_, new_n266_, new_n5690_, new_n544_, new_n4242_, new_n472_, new_n2688_, new_n5921_, y[1], new_n1090_, new_n1265_, new_n6152_, new_n6217_, new_n270_, new_n650_, new_n1193_, new_n877_, new_n1205_, new_n208_, new_n5779_, new_n235_, new_n3296_, new_n456_, new_n538_, new_n313_, new_n5584_, new_n196_, new_n535_, new_n285_, new_n5378_, new_n732_, new_n2126_, new_n388_, new_n4199_, new_n346_, new_n593_, new_n134_, new_n6062_, new_n224_, new_n5931_, new_n526_, new_n3530_, new_n3442_, new_n281_, new_n1301_, new_n855_, new_n5631_, new_n278_, new_n985_, new_n312_, new_n1092_, new_n303_, new_n525_, new_n188_, new_n5278_, new_n193_, new_n1038_, new_n637_, new_n4699_, new_n160_, new_n5186_, new_n173_, new_n4499_, new_n205_, new_n5796_, new_n696_, new_n3171_, new_n404_, new_n1386_, new_n222_, new_n948_, new_n157_, new_n5889_, new_n641_, new_n4117_, new_n170_, new_n1310_, new_n457_, new_n823_, new_n500_, new_n1123_, new_n1843_, new_n4597_, new_n161_, new_n5347_, new_n933_, new_n1140_, new_n189_, new_n1760_, new_n1379_, new_n2017_, new_n322_, new_n365_, new_n2172_, new_n414_, new_n1165_, new_n129_, new_n5621_, new_n123_, new_n4400_, new_n331_, new_n3747_, new_n213_, new_n2334_, v[1], new_n4606_, new_n426_, new_n4057_, new_n184_, new_n1143_, new_n1354_, new_n3258_, new_n217_, new_n1895_, new_n1624_, new_n3161_, v[0], new_n4248_, new_n300_, new_n818_, new_n89_, new_n754_, new_n984_, new_n3966_, new_n602_, new_n1700_, new_n438_, new_n692_, new_n424_, new_n4389_, new_n272_, new_n4464_, new_n88_, new_n2733_, new_n324_, new_n623_, new_n336_, new_n1019_, new_n145_, new_n5554_, new_n239_, new_n5349_, new_n1567_, new_n3482_, new_n1042_, new_n1455_, new_n245_, new_n3960_, new_n190_, new_n5813_, new_n202_, new_n5078_, new_n428_, new_n1621_, new_n467_, new_n3575_, new_n869_, new_n4717_, new_n144_, new_n1616_, new_n301_, new_n3761_, new_n263_, new_n5169_, new_n679_, new_n5534_, new_n204_, new_n4888_, new_n289_, new_n1619_, new_n187_, new_n5536_, new_n254_, new_n4369_, new_n450_, new_n932_, new_n1087_, new_n1110_, new_n1166_, new_n3590_, new_n199_, new_n545_})
387'b10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[24] = 1'b0;
387'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[24] = 1'b0;
387'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[24] = 1'b0;
default : coef[24] = 1'b1;
endcase
casez ({new_n221_, new_n1340_, new_n734_, new_n1752_, new_n267_, new_n5098_, new_n706_, new_n2649_, new_n194_, new_n2143_, new_n822_, new_n4340_, new_n225_, new_n1121_, new_n234_, new_n3348_, new_n247_, new_n737_, new_n320_, new_n4276_, new_n287_, new_n5363_, new_n1462_, new_n2964_, new_n721_, new_n2935_, new_n597_, new_n4885_, new_n455_, new_n1960_, new_n94_, new_n5021_, new_n382_, new_n4483_, new_n448_, new_n4599_, new_n1186_, new_n3353_, y[1], new_n4587_, new_n215_, new_n4017_, new_n499_, new_n1735_, new_n562_, new_n2509_, new_n331_, new_n2741_, new_n299_, new_n6198_, new_n5923_, new_n481_, new_n517_, new_n260_, new_n1729_, new_n257_, new_n1483_, u[2], new_n2800_, new_n979_, new_n1568_, new_n383_, new_n1228_, new_n275_, new_n4288_, new_n949_, new_n3051_, new_n150_, new_n1377_, new_n898_, new_n2919_, new_n1871_, new_n1922_, new_n494_, new_n1159_, new_n295_, new_n1581_, new_n1034_, new_n4186_, new_n389_, new_n1156_, new_n335_, new_n473_, new_n429_, new_n633_, new_n601_, new_n783_, new_n127_, new_n5604_, new_n616_, new_n1936_, new_n648_, new_n1040_, new_n244_, new_n5469_, new_n5445_, new_n447_, new_n1389_, new_n1103_, new_n1160_, new_n353_, new_n1647_, new_n148_, new_n2807_, new_n115_, new_n1065_, y[2], new_n377_, new_n1094_, new_n95_, new_n2560_, new_n290_, new_n2767_, new_n554_, new_n4731_, new_n505_, new_n3744_, new_n81_, new_n4620_, new_n86_, new_n4398_, new_n168_, new_n4082_, new_n171_, new_n870_, new_n5433_, new_n6286_, new_n509_, new_n3095_, new_n798_, new_n4274_, new_n373_, new_n3745_, new_n456_, new_n4419_, new_n305_, new_n5161_, new_n313_, new_n1147_, new_n445_, new_n755_, new_n5442_, new_n284_, new_n580_, new_n160_, new_n4155_, new_n113_, new_n891_, new_n565_, new_n2949_, new_n103_, new_n5853_, new_n230_, new_n626_, new_n166_, new_n5162_, new_n6044_, new_n6256_, new_n164_, new_n5873_, new_n172_, new_n1218_, new_n2889_, new_n1493_, new_n140_, new_n1826_, new_n269_, new_n414_, new_n87_, new_n6124_, new_n6153_, new_n536_, new_n2106_, new_n2903_, new_n485_, new_n2763_, new_n226_, new_n1906_, new_n342_, new_n1050_, new_n618_, new_n682_, new_n218_, new_n592_, new_n161_, new_n4818_, new_n2906_, new_n307_, new_n6134_, new_n151_, new_n547_, new_n238_, new_n772_, new_n199_, new_n5685_, new_n266_, new_n6169_, new_n261_, new_n2613_, new_n969_, new_n2734_, new_n739_, new_n4109_, new_n279_, new_n3083_, new_n306_, new_n5364_, new_n285_, new_n1900_, new_n323_, new_n4720_, new_n89_, new_n3525_, new_n656_, new_n3486_, new_n311_, new_n1401_, new_n391_, new_n2726_, new_n676_, new_n4958_, new_n312_, new_n2760_, new_n399_, new_n1162_, new_n408_, new_n3601_, new_n355_, new_n4550_, new_n175_, new_n3988_, new_n607_, new_n1648_, new_n163_, new_n612_, new_n155_, new_n4737_, new_n623_, new_n3816_, new_n280_, new_n4118_, new_n637_, new_n2592_, new_n219_, new_n4148_, new_n811_, new_n4579_, new_n457_, new_n4041_, new_n145_, new_n5401_, new_n291_, new_n2979_, new_n6258_, new_n158_, new_n5284_, new_n236_, new_n1409_, new_n246_, new_n5380_, new_n189_, new_n1113_, new_n541_, new_n3433_, new_n273_, new_n1485_, new_n359_, new_n974_, new_n278_, new_n1759_, new_n242_, new_n2720_, new_n1575_, new_n3447_, new_n217_, new_n1383_, new_n178_, new_n4592_, new_n729_, new_n1880_, new_n556_, new_n1250_, new_n467_, new_n496_, new_n123_, new_n1905_, new_n229_, new_n3383_, new_n504_, new_n1851_, new_n213_, new_n900_, new_n501_, new_n3503_, new_n364_, new_n402_, new_n325_, new_n751_, new_n149_, new_n545_, new_n190_, new_n1638_, new_n292_, new_n3133_, new_n2909_, new_n192_, new_n2733_, new_n185_, new_n233_, new_n792_, new_n1447_, new_n2611_, new_n3733_, new_n222_, new_n1676_, new_n174_, new_n5625_, new_n934_, new_n4743_, new_n471_, new_n3064_, new_n304_, new_n384_, new_n289_, new_n5050_, new_n2910_, new_n259_, new_n571_, new_n347_, new_n1082_, new_n410_, new_n2516_, new_n450_, new_n873_, new_n263_, new_n2125_, new_n204_, new_n464_, new_n333_, new_n862_, new_n237_, new_n5876_, new_n254_, new_n700_, new_n336_, new_n686_, new_n201_, new_n2587_, new_n182_, new_n3661_, new_n216_, new_n3063_, new_n629_, new_n2681_, new_n272_, new_n968_, new_n6055_, new_n346_, new_n596_, new_n187_, new_n4820_, new_n173_, new_n5412_, new_n424_, new_n533_, new_n129_, new_n4819_, new_n211_, new_n1849_, new_n527_, new_n3568_})
371'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00???????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????? : coef[25] = 1'b0;
371'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????? : coef[25] = 1'b0;
371'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???? : coef[25] = 1'b0;
371'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[25] = 1'b0;
371'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[25] = 1'b0;
default : coef[25] = 1'b1;
endcase
casez ({new_n327_, new_n4228_, new_n225_, new_n5991_, new_n635_, new_n5180_, new_n177_, new_n4890_, new_n437_, new_n2715_, new_n176_, new_n547_, new_n752_, new_n810_, new_n581_, new_n653_, new_n286_, new_n462_, new_n140_, new_n2607_, new_n179_, new_n5543_, new_n279_, new_n2148_, new_n418_, new_n4263_, new_n168_, new_n5514_, new_n106_, new_n4322_, new_n265_, new_n2106_, new_n197_, new_n1224_, new_n103_, new_n651_, new_n139_, new_n1282_, new_n86_, new_n617_, new_n428_, new_n3570_, new_n992_, new_n2710_, new_n289_, new_n5042_, new_n212_, new_n2608_, new_n734_, new_n2317_, new_n6187_, new_n166_, new_n5768_, new_n529_, new_n1636_, new_n356_, new_n746_, new_n500_, new_n948_, new_n557_, new_n2049_, new_n190_, new_n4933_, new_n123_, new_n415_, new_n178_, new_n4394_, new_n355_, new_n5047_, new_n157_, new_n5280_, new_n80_, new_n284_, new_n1378_, new_n450_, new_n497_, new_n169_, new_n1592_, new_n1605_, new_n1946_, new_n715_, new_n1393_, new_n249_, new_n1736_, new_n1250_, new_n3491_, new_n1748_, new_n2946_, new_n673_, new_n1637_, new_n160_, new_n1924_, new_n170_, new_n5160_, new_n6238_, new_n121_, new_n5869_, new_n150_, new_n4417_, new_n1805_, new_n3853_, new_n131_, new_n191_, new_n522_, new_n2314_, new_n423_, new_n3381_, new_n215_, new_n1044_, new_n597_, new_n2144_, new_n403_, new_n787_, new_n412_, new_n4303_, new_n94_, new_n506_, v[2], new_n248_, new_n1171_, new_n309_, new_n2791_, new_n6152_, new_n83_, new_n92_, new_n1058_, new_n171_, new_n6014_, new_n174_, new_n5734_, new_n226_, new_n2847_, new_n765_, new_n3980_, new_n6211_, new_n137_, new_n1754_, new_n172_, new_n699_, new_n277_, new_n1503_, new_n149_, new_n4435_, new_n184_, new_n5518_, new_n361_, new_n5400_, new_n276_, new_n1294_, new_n478_, new_n1022_, new_n145_, new_n5894_, new_n457_, new_n793_, new_n245_, new_n5783_, new_n5958_, new_n283_, new_n2237_, new_n721_, new_n1940_, new_n161_, new_n4381_, new_n159_, new_n2667_, new_n213_, new_n3900_, new_n84_, new_n189_, new_n1187_, new_n396_, new_n502_, v[1], new_n4611_, new_n318_, new_n5045_, new_n811_, new_n3288_, new_n173_, new_n5290_, new_n155_, new_n544_, new_n280_, new_n5770_, new_n95_, new_n1621_, new_n262_, new_n5777_, new_n167_, new_n2778_, new_n127_, new_n3943_, new_n1726_, new_n3299_, new_n442_, new_n716_, new_n82_, new_n183_, new_n1643_, new_n388_, new_n2139_, new_n447_, new_n1046_, new_n1871_, new_n3534_, new_n216_, new_n4732_, new_n494_, new_n1807_, new_n2482_, new_n6184_, new_n2171_, new_n481_, new_n3041_, new_n254_, new_n1358_, u[1], new_n93_, new_n898_, new_n162_, new_n1670_, new_n148_, new_n3660_, new_n353_, new_n451_, new_n290_, new_n5746_, new_n2800_, new_n815_, new_n1568_, new_n214_, new_n5725_, new_n783_, new_n1473_, new_n1867_, new_n1942_, new_n1222_, new_n2973_, new_n604_, new_n1219_, new_n489_, new_n1470_, new_n4628_, new_n85_, new_n4557_, new_n271_, new_n3600_, new_n1731_, new_n2955_, new_n454_, new_n5294_, new_n134_, new_n5198_, new_n346_, new_n978_, new_n5438_, new_n132_, new_n1560_, new_n164_, new_n2629_, new_n208_, new_n4147_, new_n89_, new_n5871_, new_n1045_, new_n3163_, new_n582_, new_n1983_, new_n270_, new_n4042_, new_n347_, new_n5529_, new_n201_, new_n866_, new_n385_, new_n6201_, new_n263_, new_n5967_, new_n204_, new_n3137_, new_n90_, new_n4079_, new_n272_, new_n323_, new_n129_, new_n2848_, new_n6055_, new_n259_, new_n1911_, new_n6246_, new_n240_, new_n3500_, new_n205_, new_n5658_, new_n253_, new_n4555_, new_n332_, new_n2670_, new_n246_, new_n6067_, new_n315_, new_n590_, new_n334_, new_n1625_, new_n144_, new_n5396_, new_n636_, new_n1125_, new_n237_, new_n1146_, new_n1000_, new_n2721_, new_n424_, new_n1053_, new_n115_, new_n3682_, new_n200_, new_n1327_, new_n118_, new_n1714_, new_n749_, new_n3496_, new_n924_, new_n1490_, new_n344_, new_n5849_, new_n6283_, new_n88_, new_n5699_, new_n1038_, new_n1566_, new_n554_, new_n1087_, new_n239_, new_n2559_, new_n258_, new_n482_})
338'b10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????110??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[26] = 1'b1;
338'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????? : coef[26] = 1'b1;
338'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[26] = 1'b1;
338'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?? : coef[26] = 1'b1;
338'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[26] = 1'b1;
default : coef[26] = 1'b0;
endcase
casez ({new_n341_, new_n2713_, new_n874_, new_n3291_, new_n88_, new_n220_, new_n494_, new_n178_, new_n5767_, new_n299_, new_n2814_, new_n118_, new_n5463_, new_n247_, new_n1351_, new_n142_, new_n4498_, new_n262_, new_n5056_, new_n225_, new_n2062_, new_n4596_, v[2], new_n99_, new_n2850_, new_n244_, new_n5763_, new_n82_, new_n614_, new_n426_, new_n4150_, new_n276_, new_n405_, new_n216_, new_n649_, new_n1873_, new_n3028_, new_n487_, new_n5729_, new_n796_, new_n1600_, new_n267_, new_n900_, new_n327_, new_n4834_, new_n496_, new_n1622_, new_n248_, new_n942_, new_n249_, new_n1154_, new_n101_, new_n121_, new_n455_, new_n1103_, new_n5120_, new_n578_, new_n1047_, new_n127_, new_n1021_, new_n287_, new_n1725_, new_n481_, new_n3872_, new_n377_, new_n1957_, new_n98_, new_n5016_, new_n308_, new_n1883_, new_n162_, new_n2136_, new_n115_, new_n5750_, new_n153_, new_n4758_, new_n316_, new_n1712_, new_n198_, new_n1483_, new_n271_, new_n4424_, new_n473_, new_n4193_, new_n505_, new_n4432_, new_n257_, new_n1729_, new_n353_, new_n952_, new_n579_, new_n1581_, new_n616_, new_n3554_, new_n339_, new_n451_, new_n488_, new_n2829_, new_n6188_, new_n388_, new_n3852_, new_n671_, new_n744_, new_n783_, new_n4589_, new_n330_, new_n769_, new_n695_, new_n2795_, x[2], new_n96_, new_n521_, new_n179_, new_n6206_, new_n284_, new_n468_, new_n168_, new_n5487_, new_n497_, new_n1158_, new_n132_, new_n5292_, new_n134_, new_n3889_, new_n177_, new_n2153_, new_n171_, new_n6011_, new_n6271_, new_n261_, new_n4427_, new_n530_, new_n1505_, new_n547_, new_n1101_, new_n2313_, new_n1200_, new_n3226_, new_n2901_, new_n285_, new_n4938_, new_n170_, new_n843_, new_n1578_, new_n2714_, new_n6208_, new_n384_, new_n445_, new_n498_, new_n1102_, new_n184_, new_n902_, new_n89_, new_n1464_, new_n375_, new_n1362_, new_n376_, new_n538_, new_n164_, new_n5002_, new_n226_, new_n1216_, new_n137_, new_n4518_, new_n266_, new_n3730_, new_n151_, new_n909_, new_n270_, new_n3182_, new_n301_, new_n848_, new_n2409_, new_n772_, new_n1134_, new_n368_, new_n5426_, new_n875_, new_n1373_, new_n140_, new_n1743_, new_n312_, new_n4504_, new_n379_, new_n1536_, new_n278_, new_n1741_, u[1], new_n2335_, new_n104_, new_n3740_, new_n6289_, new_n871_, new_n1379_, new_n190_, new_n1121_, new_n166_, new_n840_, new_n1378_, new_n2712_, new_n736_, new_n242_, new_n513_, new_n325_, new_n3545_, new_n363_, new_n2574_, new_n212_, new_n746_, new_n408_, new_n750_, new_n139_, new_n1210_, new_n223_, new_n1874_, new_n158_, new_n1448_, new_n625_, new_n1264_, new_n604_, new_n3433_, new_n511_, new_n974_, new_n245_, new_n1644_, new_n175_, new_n5562_, new_n259_, new_n4712_, new_n157_, new_n1576_, new_n265_, new_n4686_, new_n148_, new_n3247_, new_n318_, new_n6006_, new_n1629_, new_n2014_, new_n448_, new_n1757_, new_n253_, new_n4359_, new_n173_, new_n5801_, new_n159_, new_n5660_, new_n161_, new_n2806_, new_n370_, new_n1120_, new_n239_, new_n4294_, new_n396_, new_n410_, new_n210_, new_n5986_, new_n3603_, new_n202_, new_n989_, new_n155_, new_n5288_, new_n240_, new_n2687_, new_n84_, new_n255_, new_n292_, new_n222_, new_n756_, new_n532_, new_n2243_, new_n463_, new_n2944_, new_n340_, new_n3294_, new_n321_, new_n1476_, new_n205_, new_n5252_, new_n174_, new_n1221_, new_n333_, new_n2075_, new_n556_, new_n1031_, new_n189_, new_n689_, new_n272_, new_n2516_, new_n323_, new_n467_, new_n6270_, new_n246_, new_n1145_, new_n291_, new_n2520_, new_n424_, new_n1161_, new_n1950_, new_n2635_, new_n6280_, new_n167_, new_n4528_, new_n144_, new_n3724_, new_n478_, new_n1155_, new_n2910_, new_n557_, new_n3817_, new_n224_, new_n5286_, new_n303_, new_n1110_, new_n794_, new_n4880_, new_n199_, new_n3502_})
318'b11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????011??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????000????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????111???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????001?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011??????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00??????????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0?????????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????? : coef[27] = 1'b1;
318'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????? : coef[27] = 1'b1;
318'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[27] = 1'b1;
318'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[27] = 1'b1;
318'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[27] = 1'b1;
default : coef[27] = 1'b0;
endcase
casez ({new_n262_, new_n4836_, new_n648_, new_n3066_, new_n221_, new_n944_, new_n796_, new_n1068_, new_n1811_, new_n5103_, new_n223_, new_n4385_, new_n219_, new_n2802_, new_n118_, new_n4460_, new_n387_, new_n2755_, new_n2434_, new_n4596_, new_n748_, new_n4487_, new_n81_, new_n614_, new_n506_, new_n829_, new_n207_, new_n4996_, new_n267_, new_n5558_, new_n191_, new_n3362_, new_n404_, new_n632_, new_n139_, new_n1376_, new_n437_, new_n2641_, new_n6276_, new_n430_, new_n6022_, new_n712_, new_n1716_, new_n372_, new_n4194_, new_n976_, new_n1643_, new_n483_, new_n3176_, new_n142_, new_n3909_, new_n116_, new_n2146_, new_n382_, new_n4260_, new_n243_, new_n1073_, new_n339_, new_n1179_, new_n377_, new_n3723_, new_n868_, new_n3622_, new_n453_, new_n1389_, new_n757_, new_n2980_, new_n953_, new_n1952_, new_n122_, new_n2816_, new_n2510_, new_n3811_, new_n309_, new_n1150_, new_n310_, new_n378_, new_n316_, new_n725_, new_n356_, new_n2136_, new_n1976_, new_n104_, new_n3944_, v[2], new_n150_, new_n741_, new_n115_, new_n5906_, new_n679_, new_n821_, u[1], new_n3758_, new_n578_, new_n1181_, new_n169_, new_n5265_, new_n321_, new_n1157_, new_n214_, new_n4944_, new_n2440_, new_n227_, new_n1743_, new_n856_, new_n3676_, new_n638_, new_n1580_, new_n89_, new_n6126_, new_n340_, new_n5827_, new_n505_, new_n1557_, new_n148_, new_n5022_, new_n162_, new_n3715_, new_n388_, new_n1360_, new_n94_, new_n2825_, new_n1941_, new_n3335_, new_n640_, new_n1267_, new_n179_, new_n5861_, new_n269_, new_n2090_, new_n581_, new_n4510_, v[1], new_n261_, new_n525_, new_n140_, new_n5409_, new_n176_, new_n1556_, new_n760_, new_n1818_, new_n226_, new_n2095_, new_n218_, new_n335_, new_n1248_, new_n85_, new_n626_, new_n1051_, new_n3088_, new_n249_, new_n724_, new_n295_, new_n5812_, new_n266_, new_n540_, new_n164_, new_n5356_, new_n306_, new_n644_, new_n170_, new_n5952_, new_n370_, new_n521_, new_n270_, new_n2260_, new_n313_, new_n546_, new_n445_, new_n762_, new_n285_, new_n699_, new_n368_, new_n5697_, new_n6255_, new_n6233_, new_n215_, new_n1199_, new_n373_, new_n4728_, new_n113_, new_n6004_, new_n211_, new_n3065_, new_n231_, new_n4662_, new_n334_, new_n375_, new_n131_, new_n5105_, new_n311_, new_n336_, new_n484_, new_n554_, new_n1095_, new_n2575_, new_n307_, new_n1325_, new_n346_, new_n6085_, new_n151_, new_n1220_, new_n6234_, new_n182_, new_n832_, new_n204_, new_n902_, new_n455_, new_n1652_, new_n258_, new_n642_, new_n199_, new_n4429_, new_n279_, new_n1069_, new_n342_, new_n2140_, new_n88_, new_n3770_, new_n399_, new_n2508_, new_n584_, new_n4160_, new_n6251_, new_n284_, new_n895_, new_n6240_, new_n326_, new_n1092_, new_n1466_, new_n3254_, new_n230_, new_n903_, new_n166_, new_n1914_, new_n272_, new_n996_, new_n1379_, new_n2956_, new_n129_, new_n3448_, new_n160_, new_n4812_, new_n457_, new_n1637_, new_n177_, new_n4521_, new_n124_, new_n2775_, new_n564_, new_n4947_, new_n158_, new_n510_, new_n205_, new_n1672_, new_n2249_, new_n236_, new_n534_, new_n607_, new_n5273_, new_n157_, new_n670_, new_n508_, new_n1559_, new_n178_, new_n6121_, new_n144_, new_n6018_, new_n123_, new_n477_, new_n302_, new_n3232_, new_n161_, new_n5507_, new_n297_, new_n5904_, new_n5452_, new_n419_, new_n998_, new_n283_, new_n1605_, new_n2872_, new_n239_, new_n756_, new_n277_, new_n4058_, new_n217_, new_n5062_, new_n173_, new_n5618_, new_n185_, new_n365_, new_n472_, new_n717_, new_n478_, new_n5567_, new_n174_, new_n2750_, new_n268_, new_n5122_, new_n155_, new_n5980_, new_n5440_, new_n84_, new_n213_, new_n556_, new_n248_, new_n3359_, new_n202_, new_n454_, new_n300_, new_n5225_, new_n450_, new_n1999_, new_n208_, new_n738_, new_n722_, new_n1850_, new_n324_, new_n701_, new_n175_, new_n5589_, new_n420_, new_n2703_, new_n167_, new_n1912_, new_n253_, new_n4152_, new_n312_, new_n3979_, new_n145_, new_n5519_, new_n245_, new_n2762_, new_n344_, new_n5830_, new_n458_, new_n2765_, new_n241_, new_n2788_, new_n187_, new_n4002_, new_n467_, new_n4410_, new_n254_, new_n5870_, new_n238_, new_n325_, new_n641_, new_n794_, new_n222_, new_n1745_})
352'b11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????00?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????111????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????00????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? : coef[28] = 1'b1;
352'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011?????????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[28] = 1'b1;
352'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?? : coef[28] = 1'b1;
352'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[28] = 1'b1;
default : coef[28] = 1'b0;
endcase
casez ({new_n281_, new_n1030_, new_n230_, new_n3454_, new_n581_, new_n3539_, new_n228_, new_n1865_, new_n177_, new_n6108_, new_n142_, new_n2758_, new_n160_, new_n3919_, new_n1118_, new_n2504_, new_n207_, new_n3829_, new_n88_, new_n3685_, new_n1758_, new_n3353_, new_n6274_, new_n94_, new_n5233_, new_n940_, new_n4926_, new_n164_, new_n5933_, new_n552_, new_n5955_, new_n311_, new_n4456_, new_n137_, new_n5572_, new_n269_, new_n497_, new_n197_, new_n703_, new_n390_, new_n653_, new_n203_, new_n485_, new_n171_, new_n4280_, new_n1101_, new_n1355_, new_n866_, new_n1264_, new_n2528_, new_n3476_, new_n445_, new_n2059_, new_n113_, new_n624_, new_n132_, new_n5551_, new_n284_, new_n4852_, new_n189_, new_n4158_, new_n467_, new_n1092_, new_n734_, new_n4810_, new_n811_, new_n1818_, new_n773_, new_n3205_, new_n166_, new_n5728_, new_n928_, new_n1143_, new_n157_, new_n3670_, new_n186_, new_n2619_, new_n534_, new_n1637_, new_n607_, new_n2835_, new_n500_, new_n1147_, new_n1166_, new_n3579_, new_n2549_, new_n3556_, new_n364_, new_n817_, new_n408_, new_n961_, new_n425_, new_n797_, new_n236_, new_n2599_, new_n170_, new_n1899_, new_n243_, new_n5237_, new_n396_, new_n5945_, new_n163_, new_n2146_, new_n1952_, new_n2582_, new_n320_, new_n3052_, new_n387_, new_n1402_, new_n221_, new_n5837_, new_n283_, new_n2921_, new_n645_, new_n2505_, v[1], new_n4609_, new_n498_, new_n1429_, new_n367_, new_n1093_, new_n247_, new_n6137_, new_n262_, new_n1254_, new_n6284_, new_n6259_, new_n1715_, new_n3248_, new_n494_, new_n3796_, new_n194_, new_n4130_, new_n748_, new_n5319_, new_n121_, new_n3809_, new_n220_, new_n5006_, new_n227_, new_n5502_, new_n161_, new_n1786_, new_n226_, new_n5911_, new_n368_, new_n1412_, new_n376_, new_n4361_, new_n476_, new_n3824_, new_n192_, new_n5559_, new_n2896_, new_n731_, new_n6153_, new_n285_, new_n419_, new_n427_, new_n562_, new_n81_, new_n100_, new_n1495_, new_n216_, new_n1058_, new_n1158_, new_n1504_, new_n155_, new_n2028_, new_n291_, new_n501_, new_n159_, new_n1083_, new_n2542_, new_n3523_, new_n370_, new_n4252_, new_n478_, new_n5563_, new_n253_, new_n1167_, new_n350_, new_n354_, new_n1096_, new_n2642_, new_n420_, new_n3533_, y[2], new_n5275_, new_n276_, new_n5727_, new_n407_, new_n2743_, new_n2099_, new_n200_, new_n5482_, new_n271_, new_n3576_, new_n953_, new_n957_, new_n84_, new_n4767_, x[2], new_n264_, new_n381_, new_n299_, new_n1616_, new_n1871_, new_n2739_, new_n388_, new_n5423_, new_n150_, new_n1213_, new_n2440_, new_n360_, new_n4843_, new_n127_, new_n4207_, new_n2858_, new_n356_, new_n1953_, new_n162_, new_n1725_, new_n809_, new_n3164_, new_n524_, new_n527_, new_n604_, new_n5712_, new_n1382_, new_n3777_, new_n807_, new_n4330_, new_n2246_, new_n86_, new_n757_, new_n241_, new_n1670_, new_n290_, new_n2593_, new_n798_, new_n1159_, new_n82_, new_n4800_, new_n2149_, new_n148_, new_n601_, new_n118_, new_n1489_, new_n606_, new_n3581_, new_n633_, new_n769_, new_n201_, new_n5761_, new_n306_, new_n5804_, new_n140_, new_n3332_, new_n600_, new_n3084_, new_n4638_, new_n168_, new_n5628_, new_n386_, new_n4902_, new_n198_, new_n3372_, new_n134_, new_n4887_, new_n2937_, new_n4613_, new_n1069_, new_n3219_, new_n224_, new_n2828_, new_n153_, new_n1204_, new_n502_, new_n795_, new_n672_, new_n1042_, new_n433_, new_n1364_, new_n4665_, new_n246_, new_n939_, new_n208_, new_n4666_, new_n300_, new_n903_, new_n263_, new_n4206_, new_n323_, new_n5956_, new_n878_, new_n2929_, new_n89_, new_n1080_, new_n625_, new_n2930_, new_n355_, new_n3642_, new_n213_, new_n4131_, new_n190_, new_n5782_, new_n303_, new_n716_, new_n217_, new_n1348_, new_n123_, new_n4783_, new_n237_, new_n5196_, new_n144_, new_n5987_, new_n182_, new_n5067_, new_n707_, new_n1900_, new_n450_, new_n676_, new_n175_, new_n3605_, new_n326_, new_n5757_, new_n715_, new_n5322_, new_n316_, new_n2135_, new_n673_, new_n1398_, new_n258_, new_n1914_, new_n794_, new_n4102_, new_n435_, new_n4198_, new_n187_, new_n6061_, new_n199_, new_n589_})
343'b11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????10????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????01????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????0??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????011???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????111?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01??????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10??????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10????????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11????????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11??????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????01?????????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10???????????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11?????????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???????? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?????? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11???? : coef[29] = 1'b1;
343'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10?? : coef[29] = 1'b1;
343'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????11 : coef[29] = 1'b1;
default : coef[29] = 1'b0;
endcase
casez ({new_n6295_})
1'b0 : coef[30] = 1'b1;
default : coef[30] = 1'b0;
endcase
casez ({new_n6295_})
1'b0 : coef[31] = 1'b1;
default : coef[31] = 1'b0;
endcase
casez ({new_n81_, new_n95_})
2'b1? : new_n77_ = 1'b1;
2'b?1 : new_n77_ = 1'b1;
default : new_n77_ = 1'b0;
endcase
casez ({new_n486_, new_n437_})
2'b1? : new_n78_ = 1'b1;
2'b?1 : new_n78_ = 1'b1;
default : new_n78_ = 1'b0;
endcase
casez ({x[1], u[2]})
2'b11 : new_n79_ = 1'b1;
default : new_n79_ = 1'b0;
endcase
casez ({x[1], u[2]})
2'b01 : new_n80_ = 1'b1;
default : new_n80_ = 1'b0;
endcase
casez ({y[1], v[2]})
2'b11 : new_n81_ = 1'b1;
default : new_n81_ = 1'b0;
endcase
casez ({y[1], v[2]})
2'b01 : new_n82_ = 1'b1;
default : new_n82_ = 1'b0;
endcase
casez ({y[2], v[1]})
2'b11 : new_n83_ = 1'b1;
default : new_n83_ = 1'b0;
endcase
casez ({y[2], v[1]})
2'b01 : new_n84_ = 1'b1;
default : new_n84_ = 1'b0;
endcase
casez ({x[2], u[1]})
2'b11 : new_n85_ = 1'b1;
default : new_n85_ = 1'b0;
endcase
casez ({x[2], u[1]})
2'b01 : new_n86_ = 1'b1;
default : new_n86_ = 1'b0;
endcase
casez ({x[0], u[2], new_n93_})
3'b11? : new_n87_ = 1'b1;
3'b??1 : new_n87_ = 1'b1;
default : new_n87_ = 1'b0;
endcase
casez ({x[0], u[0]})
2'b11 : new_n88_ = 1'b1;
default : new_n88_ = 1'b0;
endcase
casez ({x[0], u[0]})
2'b01 : new_n89_ = 1'b1;
default : new_n89_ = 1'b0;
endcase
casez ({y[0], v[0]})
2'b11 : new_n90_ = 1'b1;
default : new_n90_ = 1'b0;
endcase
casez ({y[0], v[0]})
2'b01 : new_n91_ = 1'b1;
default : new_n91_ = 1'b0;
endcase
casez ({x[1], u[2]})
2'b00 : new_n92_ = 1'b1;
default : new_n92_ = 1'b0;
endcase
casez ({x[1], u[2]})
2'b10 : new_n93_ = 1'b1;
default : new_n93_ = 1'b0;
endcase
casez ({y[1], v[2]})
2'b10 : new_n94_ = 1'b1;
default : new_n94_ = 1'b0;
endcase
casez ({y[1], v[2]})
2'b00 : new_n95_ = 1'b1;
default : new_n95_ = 1'b0;
endcase
casez ({x[0], u[0]})
2'b00 : new_n96_ = 1'b1;
default : new_n96_ = 1'b0;
endcase
casez ({y[2], v[1]})
2'b00 : new_n97_ = 1'b1;
default : new_n97_ = 1'b0;
endcase
casez ({y[2], v[1]})
2'b10 : new_n98_ = 1'b1;
default : new_n98_ = 1'b0;
endcase
casez ({y[0], v[0]})
2'b00 : new_n99_ = 1'b1;
default : new_n99_ = 1'b0;
endcase
casez ({y[0], v[0]})
2'b10 : new_n100_ = 1'b1;
default : new_n100_ = 1'b0;
endcase
casez ({x[0], u[0]})
2'b10 : new_n101_ = 1'b1;
default : new_n101_ = 1'b0;
endcase
casez ({new_n82_, new_n84_, new_n83_, new_n94_})
4'b11?? : new_n102_ = 1'b1;
4'b??11 : new_n102_ = 1'b1;
default : new_n102_ = 1'b0;
endcase
casez ({x[2], u[1]})
2'b00 : new_n103_ = 1'b1;
default : new_n103_ = 1'b0;
endcase
casez ({x[2], u[1]})
2'b10 : new_n104_ = 1'b1;
default : new_n104_ = 1'b0;
endcase
casez ({new_n81_, new_n83_, new_n84_, new_n95_})
4'b11?? : new_n105_ = 1'b1;
4'b??11 : new_n105_ = 1'b1;
default : new_n105_ = 1'b0;
endcase
casez ({new_n231_, new_n337_})
2'b1? : new_n106_ = 1'b1;
2'b?1 : new_n106_ = 1'b1;
default : new_n106_ = 1'b0;
endcase
casez ({new_n79_, new_n92_})
2'b00 : new_n107_ = 1'b1;
default : new_n107_ = 1'b0;
endcase
casez ({x[1], new_n96_, new_n2917_})
3'b01? : new_n108_ = 1'b1;
3'b??1 : new_n108_ = 1'b1;
default : new_n108_ = 1'b0;
endcase
casez ({new_n80_, new_n93_})
2'b00 : new_n109_ = 1'b1;
default : new_n109_ = 1'b0;
endcase
casez ({new_n140_, new_n137_})
2'b1? : new_n110_ = 1'b1;
2'b?1 : new_n110_ = 1'b1;
default : new_n110_ = 1'b0;
endcase
casez ({new_n2977_, new_n2917_})
2'b1? : new_n111_ = 1'b1;
2'b?1 : new_n111_ = 1'b1;
default : new_n111_ = 1'b0;
endcase
casez ({new_n235_, new_n337_})
2'b1? : new_n112_ = 1'b1;
2'b?1 : new_n112_ = 1'b1;
default : new_n112_ = 1'b0;
endcase
casez ({new_n279_, new_n342_})
2'b1? : new_n113_ = 1'b1;
2'b?1 : new_n113_ = 1'b1;
default : new_n113_ = 1'b0;
endcase
casez ({u[0], new_n79_, u[2], new_n96_})
4'b01?? : new_n114_ = 1'b1;
4'b??01 : new_n114_ = 1'b1;
default : new_n114_ = 1'b0;
endcase
casez ({new_n79_, new_n83_})
2'b11 : new_n115_ = 1'b1;
default : new_n115_ = 1'b0;
endcase
casez ({new_n80_, new_n85_})
2'b11 : new_n116_ = 1'b1;
default : new_n116_ = 1'b0;
endcase
casez ({new_n235_, new_n106_})
2'b1? : new_n117_ = 1'b1;
2'b?1 : new_n117_ = 1'b1;
default : new_n117_ = 1'b0;
endcase
casez ({new_n79_, new_n84_})
2'b11 : new_n118_ = 1'b1;
default : new_n118_ = 1'b0;
endcase
casez ({u[1], new_n80_})
2'b01 : new_n119_ = 1'b1;
default : new_n119_ = 1'b0;
endcase
casez ({new_n91_, new_n97_})
2'b11 : new_n120_ = 1'b1;
default : new_n120_ = 1'b0;
endcase
casez ({y[1], new_n78_})
2'b00 : new_n121_ = 1'b1;
default : new_n121_ = 1'b0;
endcase
casez ({y[1], new_n78_})
2'b11 : new_n122_ = 1'b1;
default : new_n122_ = 1'b0;
endcase
casez ({new_n82_, new_n90_})
2'b11 : new_n123_ = 1'b1;
default : new_n123_ = 1'b0;
endcase
casez ({new_n81_, new_n86_})
2'b11 : new_n124_ = 1'b1;
default : new_n124_ = 1'b0;
endcase
casez ({new_n2977_, new_n108_})
2'b1? : new_n125_ = 1'b1;
2'b?1 : new_n125_ = 1'b1;
default : new_n125_ = 1'b0;
endcase
casez ({new_n85_, new_n93_})
2'b11 : new_n126_ = 1'b1;
default : new_n126_ = 1'b0;
endcase
casez ({y[0], new_n82_})
2'b11 : new_n127_ = 1'b1;
default : new_n127_ = 1'b0;
endcase
casez ({new_n91_, new_n98_})
2'b11 : new_n128_ = 1'b1;
default : new_n128_ = 1'b0;
endcase
casez ({new_n90_, new_n94_})
2'b11 : new_n129_ = 1'b1;
default : new_n129_ = 1'b0;
endcase
casez ({y[0], new_n88_})
2'b01 : new_n130_ = 1'b1;
default : new_n130_ = 1'b0;
endcase
casez ({new_n83_, new_n92_})
2'b11 : new_n131_ = 1'b1;
default : new_n131_ = 1'b0;
endcase
casez ({new_n445_, new_n285_})
2'b1? : new_n132_ = 1'b1;
2'b?1 : new_n132_ = 1'b1;
default : new_n132_ = 1'b0;
endcase
casez ({new_n84_, new_n86_})
2'b11 : new_n133_ = 1'b1;
default : new_n133_ = 1'b0;
endcase
casez ({new_n427_, new_n313_})
2'b1? : new_n134_ = 1'b1;
2'b?1 : new_n134_ = 1'b1;
default : new_n134_ = 1'b0;
endcase
casez ({x[2], new_n93_})
2'b01 : new_n135_ = 1'b1;
default : new_n135_ = 1'b0;
endcase
casez ({y[0], new_n89_})
2'b01 : new_n136_ = 1'b1;
default : new_n136_ = 1'b0;
endcase
casez ({new_n82_, new_n100_})
2'b11 : new_n137_ = 1'b1;
default : new_n137_ = 1'b0;
endcase
casez ({u[1], new_n96_})
2'b01 : new_n138_ = 1'b1;
default : new_n138_ = 1'b0;
endcase
casez ({new_n80_, new_n83_})
2'b11 : new_n139_ = 1'b1;
default : new_n139_ = 1'b0;
endcase
casez ({new_n81_, new_n99_})
2'b11 : new_n140_ = 1'b1;
default : new_n140_ = 1'b0;
endcase
casez ({y[0], new_n89_})
2'b11 : new_n141_ = 1'b1;
default : new_n141_ = 1'b0;
endcase
casez ({v[1], new_n79_})
2'b01 : new_n142_ = 1'b1;
default : new_n142_ = 1'b0;
endcase
casez ({x[2], new_n92_})
2'b11 : new_n143_ = 1'b1;
default : new_n143_ = 1'b0;
endcase
casez ({new_n81_, new_n90_})
2'b11 : new_n144_ = 1'b1;
default : new_n144_ = 1'b0;
endcase
casez ({new_n90_, new_n95_})
2'b11 : new_n145_ = 1'b1;
default : new_n145_ = 1'b0;
endcase
casez ({u[2], new_n101_})
2'b01 : new_n146_ = 1'b1;
default : new_n146_ = 1'b0;
endcase
casez ({y[0], new_n88_})
2'b11 : new_n147_ = 1'b1;
default : new_n147_ = 1'b0;
endcase
casez ({new_n79_, new_n97_})
2'b11 : new_n148_ = 1'b1;
default : new_n148_ = 1'b0;
endcase
casez ({new_n751_, new_n496_})
2'b1? : new_n149_ = 1'b1;
2'b?1 : new_n149_ = 1'b1;
default : new_n149_ = 1'b0;
endcase
casez ({new_n80_, new_n84_})
2'b11 : new_n150_ = 1'b1;
default : new_n150_ = 1'b0;
endcase
casez ({u[0], new_n104_})
2'b11 : new_n151_ = 1'b1;
default : new_n151_ = 1'b0;
endcase
casez ({x[2], new_n93_})
2'b11 : new_n152_ = 1'b1;
default : new_n152_ = 1'b0;
endcase
casez ({y[2], new_n79_})
2'b11 : new_n153_ = 1'b1;
default : new_n153_ = 1'b0;
endcase
casez ({new_n79_, new_n98_})
2'b11 : new_n154_ = 1'b1;
default : new_n154_ = 1'b0;
endcase
casez ({new_n82_, new_n91_})
2'b11 : new_n155_ = 1'b1;
default : new_n155_ = 1'b0;
endcase
casez ({new_n84_, new_n85_})
2'b11 : new_n156_ = 1'b1;
default : new_n156_ = 1'b0;
endcase
casez ({new_n77_, new_n91_})
2'b11 : new_n157_ = 1'b1;
default : new_n157_ = 1'b0;
endcase
casez ({x[0], new_n86_})
2'b01 : new_n158_ = 1'b1;
default : new_n158_ = 1'b0;
endcase
casez ({x[2], new_n96_})
2'b11 : new_n159_ = 1'b1;
default : new_n159_ = 1'b0;
endcase
casez ({x[0], new_n103_})
2'b11 : new_n160_ = 1'b1;
default : new_n160_ = 1'b0;
endcase
casez ({x[2], new_n96_})
2'b01 : new_n161_ = 1'b1;
default : new_n161_ = 1'b0;
endcase
casez ({y[2], new_n79_})
2'b01 : new_n162_ = 1'b1;
default : new_n162_ = 1'b0;
endcase
casez ({x[2], new_n92_})
2'b01 : new_n163_ = 1'b1;
default : new_n163_ = 1'b0;
endcase
casez ({v[0], new_n121_})
2'b01 : new_n164_ = 1'b1;
default : new_n164_ = 1'b0;
endcase
casez ({y[0], new_n101_})
2'b01 : new_n165_ = 1'b1;
default : new_n165_ = 1'b0;
endcase
casez ({x[0], new_n103_})
2'b01 : new_n166_ = 1'b1;
default : new_n166_ = 1'b0;
endcase
casez ({u[0], new_n103_})
2'b11 : new_n167_ = 1'b1;
default : new_n167_ = 1'b0;
endcase
casez ({v[0], new_n122_})
2'b01 : new_n168_ = 1'b1;
default : new_n168_ = 1'b0;
endcase
casez ({v[1], new_n80_})
2'b01 : new_n169_ = 1'b1;
default : new_n169_ = 1'b0;
endcase
casez ({x[0], new_n86_})
2'b11 : new_n170_ = 1'b1;
default : new_n170_ = 1'b0;
endcase
casez ({new_n77_, new_n99_})
2'b11 : new_n171_ = 1'b1;
default : new_n171_ = 1'b0;
endcase
casez ({new_n266_, new_n307_})
2'b1? : new_n172_ = 1'b1;
2'b?1 : new_n172_ = 1'b1;
default : new_n172_ = 1'b0;
endcase
casez ({new_n91_, new_n94_})
2'b11 : new_n173_ = 1'b1;
default : new_n173_ = 1'b0;
endcase
casez ({u[0], new_n85_})
2'b01 : new_n174_ = 1'b1;
default : new_n174_ = 1'b0;
endcase
casez ({new_n77_, new_n90_})
2'b01 : new_n175_ = 1'b1;
default : new_n175_ = 1'b0;
endcase
casez ({x[0], new_n104_})
2'b01 : new_n176_ = 1'b1;
default : new_n176_ = 1'b0;
endcase
casez ({x[0], new_n104_})
2'b11 : new_n177_ = 1'b1;
default : new_n177_ = 1'b0;
endcase
casez ({x[0], new_n85_})
2'b11 : new_n178_ = 1'b1;
default : new_n178_ = 1'b0;
endcase
casez ({new_n77_, new_n100_})
2'b01 : new_n179_ = 1'b1;
default : new_n179_ = 1'b0;
endcase
casez ({v[0], new_n98_})
2'b11 : new_n180_ = 1'b1;
default : new_n180_ = 1'b0;
endcase
casez ({new_n135_, new_n143_})
2'b00 : new_n181_ = 1'b1;
default : new_n181_ = 1'b0;
endcase
casez ({new_n88_, new_n104_})
2'b11 : new_n182_ = 1'b1;
default : new_n182_ = 1'b0;
endcase
casez ({new_n89_, new_n103_})
2'b11 : new_n183_ = 1'b1;
default : new_n183_ = 1'b0;
endcase
casez ({u[0], new_n86_})
2'b01 : new_n184_ = 1'b1;
default : new_n184_ = 1'b0;
endcase
casez ({new_n101_, new_n119_})
2'b11 : new_n185_ = 1'b1;
default : new_n185_ = 1'b0;
endcase
casez ({new_n77_, new_n90_})
2'b11 : new_n186_ = 1'b1;
default : new_n186_ = 1'b0;
endcase
casez ({u[0], new_n85_})
2'b11 : new_n187_ = 1'b1;
default : new_n187_ = 1'b0;
endcase
casez ({new_n1633_, new_n791_})
2'b1? : new_n188_ = 1'b1;
2'b?1 : new_n188_ = 1'b1;
default : new_n188_ = 1'b0;
endcase
casez ({new_n91_, new_n95_})
2'b11 : new_n189_ = 1'b1;
default : new_n189_ = 1'b0;
endcase
casez ({new_n81_, new_n91_})
2'b11 : new_n190_ = 1'b1;
default : new_n190_ = 1'b0;
endcase
casez ({new_n86_, new_n96_})
2'b11 : new_n191_ = 1'b1;
default : new_n191_ = 1'b0;
endcase
casez ({x[2], new_n101_})
2'b11 : new_n192_ = 1'b1;
default : new_n192_ = 1'b0;
endcase
casez ({new_n497_, new_n1039_})
2'b1? : new_n193_ = 1'b1;
2'b?1 : new_n193_ = 1'b1;
default : new_n193_ = 1'b0;
endcase
casez ({new_n80_, new_n97_})
2'b11 : new_n194_ = 1'b1;
default : new_n194_ = 1'b0;
endcase
casez ({new_n1640_, new_n501_})
2'b1? : new_n195_ = 1'b1;
2'b?1 : new_n195_ = 1'b1;
default : new_n195_ = 1'b0;
endcase
casez ({x[2], new_n88_})
2'b01 : new_n196_ = 1'b1;
default : new_n196_ = 1'b0;
endcase
casez ({new_n1637_, new_n1092_})
2'b1? : new_n197_ = 1'b1;
2'b?1 : new_n197_ = 1'b1;
default : new_n197_ = 1'b0;
endcase
casez ({u[2], new_n83_})
2'b11 : new_n198_ = 1'b1;
default : new_n198_ = 1'b0;
endcase
casez ({new_n86_, new_n88_})
2'b11 : new_n199_ = 1'b1;
default : new_n199_ = 1'b0;
endcase
casez ({x[2], new_n89_})
2'b11 : new_n200_ = 1'b1;
default : new_n200_ = 1'b0;
endcase
casez ({x[2], new_n88_})
2'b11 : new_n201_ = 1'b1;
default : new_n201_ = 1'b0;
endcase
casez ({new_n95_, new_n120_})
2'b11 : new_n202_ = 1'b1;
default : new_n202_ = 1'b0;
endcase
casez ({new_n607_, new_n556_})
2'b1? : new_n203_ = 1'b1;
2'b?1 : new_n203_ = 1'b1;
default : new_n203_ = 1'b0;
endcase
casez ({u[0], new_n86_})
2'b11 : new_n204_ = 1'b1;
default : new_n204_ = 1'b0;
endcase
casez ({v[0], new_n82_})
2'b11 : new_n205_ = 1'b1;
default : new_n205_ = 1'b0;
endcase
casez ({u[1], new_n84_})
2'b01 : new_n206_ = 1'b1;
default : new_n206_ = 1'b0;
endcase
casez ({y[2], new_n80_})
2'b01 : new_n207_ = 1'b1;
default : new_n207_ = 1'b0;
endcase
casez ({x[2], new_n89_})
2'b01 : new_n208_ = 1'b1;
default : new_n208_ = 1'b0;
endcase
casez ({u[2], new_n83_})
2'b01 : new_n209_ = 1'b1;
default : new_n209_ = 1'b0;
endcase
casez ({x[2], new_n101_})
2'b01 : new_n210_ = 1'b1;
default : new_n210_ = 1'b0;
endcase
casez ({new_n83_, new_n93_})
2'b11 : new_n211_ = 1'b1;
default : new_n211_ = 1'b0;
endcase
casez ({new_n80_, new_n98_})
2'b11 : new_n212_ = 1'b1;
default : new_n212_ = 1'b0;
endcase
casez ({v[0], new_n94_})
2'b11 : new_n213_ = 1'b1;
default : new_n213_ = 1'b0;
endcase
casez ({v[1], new_n92_})
2'b01 : new_n214_ = 1'b1;
default : new_n214_ = 1'b0;
endcase
casez ({new_n85_, new_n96_})
2'b11 : new_n215_ = 1'b1;
default : new_n215_ = 1'b0;
endcase
casez ({y[2], new_n80_})
2'b11 : new_n216_ = 1'b1;
default : new_n216_ = 1'b0;
endcase
casez ({v[0], new_n95_})
2'b11 : new_n217_ = 1'b1;
default : new_n217_ = 1'b0;
endcase
casez ({new_n95_, new_n99_})
2'b11 : new_n218_ = 1'b1;
default : new_n218_ = 1'b0;
endcase
casez ({new_n92_, new_n97_})
2'b11 : new_n219_ = 1'b1;
default : new_n219_ = 1'b0;
endcase
casez ({y[0], new_n94_})
2'b11 : new_n220_ = 1'b1;
default : new_n220_ = 1'b0;
endcase
casez ({y[0], new_n81_})
2'b01 : new_n221_ = 1'b1;
default : new_n221_ = 1'b0;
endcase
casez ({v[2], new_n90_})
2'b11 : new_n222_ = 1'b1;
default : new_n222_ = 1'b0;
endcase
casez ({x[0], new_n85_})
2'b01 : new_n223_ = 1'b1;
default : new_n223_ = 1'b0;
endcase
casez ({u[0], u[1]})
2'b11 : new_n224_ = 1'b1;
default : new_n224_ = 1'b0;
endcase
casez ({y[0], new_n77_})
2'b10 : new_n225_ = 1'b1;
default : new_n225_ = 1'b0;
endcase
casez ({new_n94_, new_n100_})
2'b11 : new_n226_ = 1'b1;
default : new_n226_ = 1'b0;
endcase
casez ({new_n486_, new_n94_})
2'b1? : new_n227_ = 1'b1;
2'b?1 : new_n227_ = 1'b1;
default : new_n227_ = 1'b0;
endcase
casez ({y[0], new_n82_})
2'b01 : new_n228_ = 1'b1;
default : new_n228_ = 1'b0;
endcase
casez ({new_n85_, new_n101_})
2'b11 : new_n229_ = 1'b1;
default : new_n229_ = 1'b0;
endcase
casez ({x[0], u[1]})
2'b00 : new_n230_ = 1'b1;
default : new_n230_ = 1'b0;
endcase
casez ({y[1], new_n99_})
2'b01 : new_n231_ = 1'b1;
default : new_n231_ = 1'b0;
endcase
casez ({new_n697_, new_n355_})
2'b1? : new_n232_ = 1'b1;
2'b?1 : new_n232_ = 1'b1;
default : new_n232_ = 1'b0;
endcase
casez ({y[2], new_n500_, new_n123_})
3'b11? : new_n233_ = 1'b1;
3'b??1 : new_n233_ = 1'b1;
default : new_n233_ = 1'b0;
endcase
casez ({u[0], u[1]})
2'b00 : new_n234_ = 1'b1;
default : new_n234_ = 1'b0;
endcase
casez ({y[1], new_n100_})
2'b11 : new_n235_ = 1'b1;
default : new_n235_ = 1'b0;
endcase
casez ({x[0], new_n126_})
2'b01 : new_n236_ = 1'b1;
default : new_n236_ = 1'b0;
endcase
casez ({new_n89_, new_n104_})
2'b11 : new_n237_ = 1'b1;
default : new_n237_ = 1'b0;
endcase
casez ({new_n85_, new_n89_})
2'b11 : new_n238_ = 1'b1;
default : new_n238_ = 1'b0;
endcase
casez ({v[0], new_n81_})
2'b11 : new_n239_ = 1'b1;
default : new_n239_ = 1'b0;
endcase
casez ({v[2], new_n90_})
2'b01 : new_n240_ = 1'b1;
default : new_n240_ = 1'b0;
endcase
casez ({y[2], new_n92_})
2'b11 : new_n241_ = 1'b1;
default : new_n241_ = 1'b0;
endcase
casez ({x[0], u[1]})
2'b10 : new_n242_ = 1'b1;
default : new_n242_ = 1'b0;
endcase
casez ({new_n84_, new_n93_})
2'b11 : new_n243_ = 1'b1;
default : new_n243_ = 1'b0;
endcase
casez ({y[0], new_n81_})
2'b11 : new_n244_ = 1'b1;
default : new_n244_ = 1'b0;
endcase
casez ({new_n98_, new_n129_})
2'b11 : new_n245_ = 1'b1;
default : new_n245_ = 1'b0;
endcase
casez ({v[0], new_n121_})
2'b11 : new_n246_ = 1'b1;
default : new_n246_ = 1'b0;
endcase
casez ({y[0], new_n95_})
2'b01 : new_n247_ = 1'b1;
default : new_n247_ = 1'b0;
endcase
casez ({new_n86_, new_n101_})
2'b11 : new_n248_ = 1'b1;
default : new_n248_ = 1'b0;
endcase
casez ({y[2], new_n92_})
2'b01 : new_n249_ = 1'b1;
default : new_n249_ = 1'b0;
endcase
casez ({v[1], new_n93_})
2'b01 : new_n250_ = 1'b1;
default : new_n250_ = 1'b0;
endcase
casez ({new_n88_, new_n103_})
2'b11 : new_n251_ = 1'b1;
default : new_n251_ = 1'b0;
endcase
casez ({new_n127_, new_n140_})
2'b00 : new_n252_ = 1'b1;
default : new_n252_ = 1'b0;
endcase
casez ({new_n81_, new_n120_})
2'b11 : new_n253_ = 1'b1;
default : new_n253_ = 1'b0;
endcase
casez ({u[1], new_n89_})
2'b11 : new_n254_ = 1'b1;
default : new_n254_ = 1'b0;
endcase
casez ({v[2], new_n91_})
2'b11 : new_n255_ = 1'b1;
default : new_n255_ = 1'b0;
endcase
casez ({new_n396_, new_n751_})
2'b1? : new_n256_ = 1'b1;
2'b?1 : new_n256_ = 1'b1;
default : new_n256_ = 1'b0;
endcase
casez ({u[2], v[1]})
2'b00 : new_n257_ = 1'b1;
default : new_n257_ = 1'b0;
endcase
casez ({u[1], new_n88_})
2'b11 : new_n258_ = 1'b1;
default : new_n258_ = 1'b0;
endcase
casez ({new_n77_, new_n120_})
2'b01 : new_n259_ = 1'b1;
default : new_n259_ = 1'b0;
endcase
casez ({u[2], v[1]})
2'b10 : new_n260_ = 1'b1;
default : new_n260_ = 1'b0;
endcase
casez ({new_n82_, new_n99_})
2'b11 : new_n261_ = 1'b1;
default : new_n261_ = 1'b0;
endcase
casez ({y[0], new_n95_})
2'b11 : new_n262_ = 1'b1;
default : new_n262_ = 1'b0;
endcase
casez ({v[0], new_n122_})
2'b11 : new_n263_ = 1'b1;
default : new_n263_ = 1'b0;
endcase
casez ({x[1], new_n83_})
2'b11 : new_n264_ = 1'b1;
default : new_n264_ = 1'b0;
endcase
casez ({x[0], new_n116_})
2'b11 : new_n265_ = 1'b1;
default : new_n265_ = 1'b0;
endcase
casez ({v[0], new_n94_})
2'b01 : new_n266_ = 1'b1;
default : new_n266_ = 1'b0;
endcase
casez ({y[0], new_n77_})
2'b01 : new_n267_ = 1'b1;
default : new_n267_ = 1'b0;
endcase
casez ({u[0], new_n126_})
2'b01 : new_n268_ = 1'b1;
default : new_n268_ = 1'b0;
endcase
casez ({new_n100_, new_n105_})
2'b11 : new_n269_ = 1'b1;
default : new_n269_ = 1'b0;
endcase
casez ({new_n99_, new_n102_})
2'b11 : new_n270_ = 1'b1;
default : new_n270_ = 1'b0;
endcase
casez ({new_n81_, new_n130_})
2'b11 : new_n271_ = 1'b1;
default : new_n271_ = 1'b0;
endcase
casez ({new_n77_, new_n128_})
2'b01 : new_n272_ = 1'b1;
default : new_n272_ = 1'b0;
endcase
casez ({v[1], new_n79_})
2'b11 : new_n273_ = 1'b1;
default : new_n273_ = 1'b0;
endcase
casez ({u[2], new_n97_})
2'b01 : new_n274_ = 1'b1;
default : new_n274_ = 1'b0;
endcase
casez ({new_n84_, new_n92_})
2'b11 : new_n275_ = 1'b1;
default : new_n275_ = 1'b0;
endcase
casez ({new_n1504_, new_n350_})
2'b1? : new_n276_ = 1'b1;
2'b?1 : new_n276_ = 1'b1;
default : new_n276_ = 1'b0;
endcase
casez ({u[1], new_n111_})
2'b01 : new_n277_ = 1'b1;
default : new_n277_ = 1'b0;
endcase
casez ({x[0], x[2]})
2'b11 : new_n278_ = 1'b1;
default : new_n278_ = 1'b0;
endcase
casez ({v[0], new_n95_})
2'b01 : new_n279_ = 1'b1;
default : new_n279_ = 1'b0;
endcase
casez ({new_n81_, new_n128_})
2'b11 : new_n280_ = 1'b1;
default : new_n280_ = 1'b0;
endcase
casez ({x[0], x[2]})
2'b00 : new_n281_ = 1'b1;
default : new_n281_ = 1'b0;
endcase
casez ({new_n83_, new_n135_})
2'b11 : new_n282_ = 1'b1;
default : new_n282_ = 1'b0;
endcase
casez ({u[1], new_n108_})
2'b01 : new_n283_ = 1'b1;
default : new_n283_ = 1'b0;
endcase
casez ({x[0], x[2]})
2'b10 : new_n284_ = 1'b1;
default : new_n284_ = 1'b0;
endcase
casez ({v[2], new_n100_})
2'b01 : new_n285_ = 1'b1;
default : new_n285_ = 1'b0;
endcase
casez ({x[0], new_n116_})
2'b01 : new_n286_ = 1'b1;
default : new_n286_ = 1'b0;
endcase
casez ({u[2], new_n97_})
2'b11 : new_n287_ = 1'b1;
default : new_n287_ = 1'b0;
endcase
casez ({new_n193_, new_n203_})
2'b00 : new_n288_ = 1'b1;
default : new_n288_ = 1'b0;
endcase
casez ({new_n98_, new_n123_})
2'b11 : new_n289_ = 1'b1;
default : new_n289_ = 1'b0;
endcase
casez ({new_n81_, new_n136_})
2'b11 : new_n290_ = 1'b1;
default : new_n290_ = 1'b0;
endcase
casez ({new_n545_, new_n325_})
2'b1? : new_n291_ = 1'b1;
2'b?1 : new_n291_ = 1'b1;
default : new_n291_ = 1'b0;
endcase
casez ({x[1], new_n138_})
2'b01 : new_n292_ = 1'b1;
default : new_n292_ = 1'b0;
endcase
casez ({new_n86_, new_n89_})
2'b11 : new_n293_ = 1'b1;
default : new_n293_ = 1'b0;
endcase
casez ({new_n99_, new_n124_})
2'b11 : new_n294_ = 1'b1;
default : new_n294_ = 1'b0;
endcase
casez ({new_n80_, new_n133_})
2'b11 : new_n295_ = 1'b1;
default : new_n295_ = 1'b0;
endcase
casez ({y[1], new_n128_, new_n1944_})
3'b11? : new_n296_ = 1'b1;
3'b??1 : new_n296_ = 1'b1;
default : new_n296_ = 1'b0;
endcase
casez ({new_n1163_, new_n536_})
2'b1? : new_n297_ = 1'b1;
2'b?1 : new_n297_ = 1'b1;
default : new_n297_ = 1'b0;
endcase
casez ({new_n1166_, new_n233_})
2'b1? : new_n298_ = 1'b1;
2'b?1 : new_n298_ = 1'b1;
default : new_n298_ = 1'b0;
endcase
casez ({y[0], new_n94_})
2'b01 : new_n299_ = 1'b1;
default : new_n299_ = 1'b0;
endcase
casez ({x[2], u[0]})
2'b01 : new_n300_ = 1'b1;
default : new_n300_ = 1'b0;
endcase
casez ({u[1], new_n89_})
2'b01 : new_n301_ = 1'b1;
default : new_n301_ = 1'b0;
endcase
casez ({new_n161_, new_n176_})
2'b00 : new_n302_ = 1'b1;
default : new_n302_ = 1'b0;
endcase
casez ({new_n82_, new_n128_})
2'b11 : new_n303_ = 1'b1;
default : new_n303_ = 1'b0;
endcase
casez ({new_n90_, new_n227_})
2'b00 : new_n304_ = 1'b1;
default : new_n304_ = 1'b0;
endcase
casez ({x[0], x[2]})
2'b01 : new_n305_ = 1'b1;
default : new_n305_ = 1'b0;
endcase
casez ({new_n81_, new_n100_})
2'b11 : new_n306_ = 1'b1;
default : new_n306_ = 1'b0;
endcase
casez ({v[2], new_n100_})
2'b11 : new_n307_ = 1'b1;
default : new_n307_ = 1'b0;
endcase
casez ({new_n103_, new_n141_})
2'b11 : new_n308_ = 1'b1;
default : new_n308_ = 1'b0;
endcase
casez ({new_n92_, new_n98_})
2'b11 : new_n309_ = 1'b1;
default : new_n309_ = 1'b0;
endcase
casez ({new_n84_, new_n119_})
2'b11 : new_n310_ = 1'b1;
default : new_n310_ = 1'b0;
endcase
casez ({v[1], new_n137_})
2'b01 : new_n311_ = 1'b1;
default : new_n311_ = 1'b0;
endcase
casez ({new_n91_, new_n102_})
2'b11 : new_n312_ = 1'b1;
default : new_n312_ = 1'b0;
endcase
casez ({v[2], new_n99_})
2'b01 : new_n313_ = 1'b1;
default : new_n313_ = 1'b0;
endcase
casez ({new_n1401_, new_n199_})
2'b1? : new_n314_ = 1'b1;
2'b?1 : new_n314_ = 1'b1;
default : new_n314_ = 1'b0;
endcase
casez ({y[1], v[0]})
2'b11 : new_n315_ = 1'b1;
default : new_n315_ = 1'b0;
endcase
casez ({u[2], new_n84_})
2'b11 : new_n316_ = 1'b1;
default : new_n316_ = 1'b0;
endcase
casez ({new_n93_, new_n97_})
2'b11 : new_n317_ = 1'b1;
default : new_n317_ = 1'b0;
endcase
casez ({v[2], new_n91_})
2'b01 : new_n318_ = 1'b1;
default : new_n318_ = 1'b0;
endcase
casez ({new_n94_, new_n127_})
2'b00 : new_n319_ = 1'b1;
default : new_n319_ = 1'b0;
endcase
casez ({new_n95_, new_n244_})
2'b00 : new_n320_ = 1'b1;
default : new_n320_ = 1'b0;
endcase
casez ({y[2], new_n93_})
2'b01 : new_n321_ = 1'b1;
default : new_n321_ = 1'b0;
endcase
casez ({new_n414_, new_n675_})
2'b1? : new_n322_ = 1'b1;
2'b?1 : new_n322_ = 1'b1;
default : new_n322_ = 1'b0;
endcase
casez ({u[0], new_n152_})
2'b11 : new_n323_ = 1'b1;
default : new_n323_ = 1'b0;
endcase
casez ({new_n88_, new_n135_})
2'b11 : new_n324_ = 1'b1;
default : new_n324_ = 1'b0;
endcase
casez ({new_n95_, new_n128_})
2'b11 : new_n325_ = 1'b1;
default : new_n325_ = 1'b0;
endcase
casez ({new_n545_, new_n289_})
2'b1? : new_n326_ = 1'b1;
2'b?1 : new_n326_ = 1'b1;
default : new_n326_ = 1'b0;
endcase
casez ({new_n648_, new_n270_})
2'b1? : new_n327_ = 1'b1;
2'b?1 : new_n327_ = 1'b1;
default : new_n327_ = 1'b0;
endcase
casez ({y[2], u[2]})
2'b11 : new_n328_ = 1'b1;
default : new_n328_ = 1'b0;
endcase
casez ({new_n104_, new_n147_})
2'b11 : new_n329_ = 1'b1;
default : new_n329_ = 1'b0;
endcase
casez ({new_n82_, new_n130_})
2'b11 : new_n330_ = 1'b1;
default : new_n330_ = 1'b0;
endcase
casez ({u[1], new_n125_})
2'b01 : new_n331_ = 1'b1;
default : new_n331_ = 1'b0;
endcase
casez ({y[2], u[2]})
2'b01 : new_n332_ = 1'b1;
default : new_n332_ = 1'b0;
endcase
casez ({new_n205_, new_n240_})
2'b00 : new_n333_ = 1'b1;
default : new_n333_ = 1'b0;
endcase
casez ({new_n89_, new_n143_})
2'b11 : new_n334_ = 1'b1;
default : new_n334_ = 1'b0;
endcase
casez ({new_n92_, new_n133_})
2'b11 : new_n335_ = 1'b1;
default : new_n335_ = 1'b0;
endcase
casez ({new_n88_, new_n143_})
2'b11 : new_n336_ = 1'b1;
default : new_n336_ = 1'b0;
endcase
casez ({v[0], v[2]})
2'b00 : new_n337_ = 1'b1;
default : new_n337_ = 1'b0;
endcase
casez ({x[1], new_n83_})
2'b01 : new_n338_ = 1'b1;
default : new_n338_ = 1'b0;
endcase
casez ({new_n82_, new_n136_})
2'b11 : new_n339_ = 1'b1;
default : new_n339_ = 1'b0;
endcase
casez ({new_n84_, new_n116_})
2'b11 : new_n340_ = 1'b1;
default : new_n340_ = 1'b0;
endcase
casez ({new_n487_, new_n82_})
2'b1? : new_n341_ = 1'b1;
2'b?1 : new_n341_ = 1'b1;
default : new_n341_ = 1'b0;
endcase
casez ({v[2], new_n99_})
2'b11 : new_n342_ = 1'b1;
default : new_n342_ = 1'b0;
endcase
casez ({new_n93_, new_n98_})
2'b11 : new_n343_ = 1'b1;
default : new_n343_ = 1'b0;
endcase
casez ({u[1], new_n88_})
2'b01 : new_n344_ = 1'b1;
default : new_n344_ = 1'b0;
endcase
casez ({new_n83_, new_n119_})
2'b11 : new_n345_ = 1'b1;
default : new_n345_ = 1'b0;
endcase
casez ({u[0], u[1]})
2'b10 : new_n346_ = 1'b1;
default : new_n346_ = 1'b0;
endcase
casez ({new_n85_, new_n88_})
2'b11 : new_n347_ = 1'b1;
default : new_n347_ = 1'b0;
endcase
casez ({new_n119_, new_n163_})
2'b00 : new_n348_ = 1'b1;
default : new_n348_ = 1'b0;
endcase
casez ({x[0], new_n109_, new_n107_})
3'b11? : new_n349_ = 1'b1;
3'b0?1 : new_n349_ = 1'b1;
default : new_n349_ = 1'b0;
endcase
casez ({new_n86_, new_n146_})
2'b11 : new_n350_ = 1'b1;
default : new_n350_ = 1'b0;
endcase
casez ({new_n522_, v[2]})
2'b1? : new_n351_ = 1'b1;
2'b?0 : new_n351_ = 1'b1;
default : new_n351_ = 1'b0;
endcase
casez ({new_n90_, new_n124_})
2'b11 : new_n352_ = 1'b1;
default : new_n352_ = 1'b0;
endcase
casez ({new_n95_, new_n136_})
2'b11 : new_n353_ = 1'b1;
default : new_n353_ = 1'b0;
endcase
casez ({new_n1605_, new_n303_})
2'b1? : new_n354_ = 1'b1;
2'b?1 : new_n354_ = 1'b1;
default : new_n354_ = 1'b0;
endcase
casez ({new_n98_, new_n186_})
2'b11 : new_n355_ = 1'b1;
default : new_n355_ = 1'b0;
endcase
casez ({y[2], new_n93_})
2'b11 : new_n356_ = 1'b1;
default : new_n356_ = 1'b0;
endcase
casez ({u[1], new_n101_})
2'b01 : new_n357_ = 1'b1;
default : new_n357_ = 1'b0;
endcase
casez ({u[2], new_n84_})
2'b01 : new_n358_ = 1'b1;
default : new_n358_ = 1'b0;
endcase
casez ({new_n213_, new_n222_})
2'b00 : new_n359_ = 1'b1;
default : new_n359_ = 1'b0;
endcase
casez ({y[0], new_n77_})
2'b11 : new_n360_ = 1'b1;
default : new_n360_ = 1'b0;
endcase
casez ({y[1], new_n180_})
2'b01 : new_n361_ = 1'b1;
default : new_n361_ = 1'b0;
endcase
casez ({x[1], y[1], new_n100_, new_n337_})
4'b001? : new_n362_ = 1'b1;
4'b???1 : new_n362_ = 1'b1;
default : new_n362_ = 1'b0;
endcase
casez ({v[1], new_n80_})
2'b11 : new_n363_ = 1'b1;
default : new_n363_ = 1'b0;
endcase
casez ({new_n217_, new_n255_})
2'b00 : new_n364_ = 1'b1;
default : new_n364_ = 1'b0;
endcase
casez ({new_n636_, new_n84_, new_n205_})
3'b1?? : new_n365_ = 1'b1;
3'b?11 : new_n365_ = 1'b1;
default : new_n365_ = 1'b0;
endcase
casez ({new_n84_, new_n135_})
2'b11 : new_n366_ = 1'b1;
default : new_n366_ = 1'b0;
endcase
casez ({new_n115_, new_n138_})
2'b11 : new_n367_ = 1'b1;
default : new_n367_ = 1'b0;
endcase
casez ({v[1], new_n110_})
2'b01 : new_n368_ = 1'b1;
default : new_n368_ = 1'b0;
endcase
casez ({x[1], new_n84_})
2'b11 : new_n369_ = 1'b1;
default : new_n369_ = 1'b0;
endcase
casez ({new_n159_, new_n166_})
2'b00 : new_n370_ = 1'b1;
default : new_n370_ = 1'b0;
endcase
casez ({new_n94_, new_n141_})
2'b11 : new_n371_ = 1'b1;
default : new_n371_ = 1'b0;
endcase
casez ({new_n82_, new_n165_})
2'b11 : new_n372_ = 1'b1;
default : new_n372_ = 1'b0;
endcase
casez ({v[1], new_n112_})
2'b01 : new_n373_ = 1'b1;
default : new_n373_ = 1'b0;
endcase
casez ({new_n115_, new_n168_, new_n118_, new_n164_})
4'b11?? : new_n374_ = 1'b1;
4'b??11 : new_n374_ = 1'b1;
default : new_n374_ = 1'b0;
endcase
casez ({v[1], new_n117_})
2'b01 : new_n375_ = 1'b1;
default : new_n375_ = 1'b0;
endcase
casez ({new_n1403_, new_n3606_})
2'b1? : new_n376_ = 1'b1;
2'b?1 : new_n376_ = 1'b1;
default : new_n376_ = 1'b0;
endcase
casez ({new_n81_, new_n141_})
2'b11 : new_n377_ = 1'b1;
default : new_n377_ = 1'b0;
endcase
casez ({new_n94_, new_n136_})
2'b11 : new_n378_ = 1'b1;
default : new_n378_ = 1'b0;
endcase
casez ({new_n674_, new_n126_})
2'b1? : new_n379_ = 1'b1;
2'b?1 : new_n379_ = 1'b1;
default : new_n379_ = 1'b0;
endcase
casez ({new_n190_, new_n217_})
2'b00 : new_n380_ = 1'b1;
default : new_n380_ = 1'b0;
endcase
casez ({new_n94_, new_n130_})
2'b11 : new_n381_ = 1'b1;
default : new_n381_ = 1'b0;
endcase
casez ({new_n83_, new_n116_})
2'b11 : new_n382_ = 1'b1;
default : new_n382_ = 1'b0;
endcase
casez ({u[2], new_n156_})
2'b11 : new_n383_ = 1'b1;
default : new_n383_ = 1'b0;
endcase
casez ({new_n118_, new_n138_})
2'b11 : new_n384_ = 1'b1;
default : new_n384_ = 1'b0;
endcase
casez ({x[2], u[0]})
2'b11 : new_n385_ = 1'b1;
default : new_n385_ = 1'b0;
endcase
casez ({new_n95_, new_n100_})
2'b11 : new_n386_ = 1'b1;
default : new_n386_ = 1'b0;
endcase
casez ({new_n81_, new_n165_})
2'b11 : new_n387_ = 1'b1;
default : new_n387_ = 1'b0;
endcase
casez ({new_n83_, new_n109_})
2'b10 : new_n388_ = 1'b1;
default : new_n388_ = 1'b0;
endcase
casez ({new_n95_, new_n130_})
2'b11 : new_n389_ = 1'b1;
default : new_n389_ = 1'b0;
endcase
casez ({u[2], new_n133_})
2'b11 : new_n390_ = 1'b1;
default : new_n390_ = 1'b0;
endcase
casez ({v[1], new_n140_})
2'b01 : new_n391_ = 1'b1;
default : new_n391_ = 1'b0;
endcase
casez ({new_n875_, new_n538_})
2'b1? : new_n392_ = 1'b1;
2'b?1 : new_n392_ = 1'b1;
default : new_n392_ = 1'b0;
endcase
casez ({new_n231_, new_n279_})
2'b00 : new_n393_ = 1'b1;
default : new_n393_ = 1'b0;
endcase
casez ({new_n144_, new_n217_})
2'b00 : new_n394_ = 1'b1;
default : new_n394_ = 1'b0;
endcase
casez ({new_n103_, new_n147_})
2'b11 : new_n395_ = 1'b1;
default : new_n395_ = 1'b0;
endcase
casez ({x[2], new_n146_})
2'b11 : new_n396_ = 1'b1;
default : new_n396_ = 1'b0;
endcase
casez ({x[0], new_n124_})
2'b11 : new_n397_ = 1'b1;
default : new_n397_ = 1'b0;
endcase
casez ({new_n83_, new_n107_})
2'b10 : new_n398_ = 1'b1;
default : new_n398_ = 1'b0;
endcase
casez ({new_n467_, new_n545_})
2'b1? : new_n399_ = 1'b1;
2'b?1 : new_n399_ = 1'b1;
default : new_n399_ = 1'b0;
endcase
casez ({new_n2154_, new_n298_})
2'b1? : new_n400_ = 1'b1;
2'b?1 : new_n400_ = 1'b1;
default : new_n400_ = 1'b0;
endcase
casez ({x[2], u[0]})
2'b00 : new_n401_ = 1'b1;
default : new_n401_ = 1'b0;
endcase
casez ({new_n1043_, new_n2687_})
2'b1? : new_n402_ = 1'b1;
2'b?1 : new_n402_ = 1'b1;
default : new_n402_ = 1'b0;
endcase
casez ({new_n504_, new_n556_})
2'b1? : new_n403_ = 1'b1;
2'b?1 : new_n403_ = 1'b1;
default : new_n403_ = 1'b0;
endcase
casez ({new_n93_, new_n133_})
2'b11 : new_n404_ = 1'b1;
default : new_n404_ = 1'b0;
endcase
casez ({new_n98_, new_n127_})
2'b11 : new_n405_ = 1'b1;
default : new_n405_ = 1'b0;
endcase
casez ({new_n288_, new_n314_})
2'b10 : new_n406_ = 1'b1;
default : new_n406_ = 1'b0;
endcase
casez ({new_n84_, new_n163_})
2'b11 : new_n407_ = 1'b1;
default : new_n407_ = 1'b0;
endcase
casez ({x[0], new_n124_})
2'b01 : new_n408_ = 1'b1;
default : new_n408_ = 1'b0;
endcase
casez ({new_n202_, new_n280_})
2'b00 : new_n409_ = 1'b1;
default : new_n409_ = 1'b0;
endcase
casez ({new_n253_, new_n312_})
2'b00 : new_n410_ = 1'b1;
default : new_n410_ = 1'b0;
endcase
casez ({y[2], u[2]})
2'b10 : new_n411_ = 1'b1;
default : new_n411_ = 1'b0;
endcase
casez ({new_n1126_, new_n1902_})
2'b1? : new_n412_ = 1'b1;
2'b?1 : new_n412_ = 1'b1;
default : new_n412_ = 1'b0;
endcase
casez ({new_n177_, new_n210_})
2'b00 : new_n413_ = 1'b1;
default : new_n413_ = 1'b0;
endcase
casez ({x[2], new_n146_})
2'b01 : new_n414_ = 1'b1;
default : new_n414_ = 1'b0;
endcase
casez ({x[0], new_n517_, new_n340_})
3'b11? : new_n415_ = 1'b1;
3'b??1 : new_n415_ = 1'b1;
default : new_n415_ = 1'b0;
endcase
casez ({y[0], new_n102_})
2'b01 : new_n416_ = 1'b1;
default : new_n416_ = 1'b0;
endcase
casez ({x[1], new_n84_})
2'b01 : new_n417_ = 1'b1;
default : new_n417_ = 1'b0;
endcase
casez ({new_n160_, new_n192_})
2'b00 : new_n418_ = 1'b1;
default : new_n418_ = 1'b0;
endcase
casez ({new_n138_, new_n162_})
2'b11 : new_n419_ = 1'b1;
default : new_n419_ = 1'b0;
endcase
casez ({new_n78_, new_n315_})
2'b01 : new_n420_ = 1'b1;
default : new_n420_ = 1'b0;
endcase
casez ({new_n96_, new_n124_})
2'b11 : new_n421_ = 1'b1;
default : new_n421_ = 1'b0;
endcase
casez ({new_n77_, new_n91_})
2'b01 : new_n422_ = 1'b1;
default : new_n422_ = 1'b0;
endcase
casez ({new_n84_, new_n126_})
2'b11 : new_n423_ = 1'b1;
default : new_n423_ = 1'b0;
endcase
casez ({new_n89_, new_n135_})
2'b11 : new_n424_ = 1'b1;
default : new_n424_ = 1'b0;
endcase
casez ({new_n984_, new_n272_})
2'b1? : new_n425_ = 1'b1;
2'b?1 : new_n425_ = 1'b1;
default : new_n425_ = 1'b0;
endcase
casez ({new_n86_, new_n114_})
2'b11 : new_n426_ = 1'b1;
default : new_n426_ = 1'b0;
endcase
casez ({v[0], new_n81_})
2'b01 : new_n427_ = 1'b1;
default : new_n427_ = 1'b0;
endcase
casez ({new_n239_, new_n240_})
2'b00 : new_n428_ = 1'b1;
default : new_n428_ = 1'b0;
endcase
casez ({new_n92_, new_n156_})
2'b11 : new_n429_ = 1'b1;
default : new_n429_ = 1'b0;
endcase
casez ({v[1], new_n109_})
2'b00 : new_n430_ = 1'b1;
default : new_n430_ = 1'b0;
endcase
casez ({new_n2934_, new_n86_})
2'b1? : new_n431_ = 1'b1;
2'b?1 : new_n431_ = 1'b1;
default : new_n431_ = 1'b0;
endcase
casez ({new_n79_, new_n83_})
2'b01 : new_n432_ = 1'b1;
default : new_n432_ = 1'b0;
endcase
casez ({new_n82_, new_n91_})
2'b01 : new_n433_ = 1'b1;
default : new_n433_ = 1'b0;
endcase
casez ({new_n2757_, new_n3592_})
2'b1? : new_n434_ = 1'b1;
2'b?1 : new_n434_ = 1'b1;
default : new_n434_ = 1'b0;
endcase
casez ({v[1], new_n116_})
2'b01 : new_n435_ = 1'b1;
default : new_n435_ = 1'b0;
endcase
casez ({u[0], u[1], new_n349_})
3'b1?? : new_n436_ = 1'b1;
3'b?10 : new_n436_ = 1'b1;
default : new_n436_ = 1'b0;
endcase
casez ({y[0], v[2]})
2'b00 : new_n437_ = 1'b1;
default : new_n437_ = 1'b0;
endcase
casez ({y[1], new_n91_})
2'b01 : new_n438_ = 1'b1;
default : new_n438_ = 1'b0;
endcase
casez ({new_n235_, new_n266_})
2'b00 : new_n439_ = 1'b1;
default : new_n439_ = 1'b0;
endcase
casez ({new_n1602_, new_n3516_})
2'b1? : new_n440_ = 1'b1;
2'b?1 : new_n440_ = 1'b1;
default : new_n440_ = 1'b0;
endcase
casez ({y[2], new_n116_})
2'b01 : new_n441_ = 1'b1;
default : new_n441_ = 1'b0;
endcase
casez ({new_n97_, new_n127_})
2'b11 : new_n442_ = 1'b1;
default : new_n442_ = 1'b0;
endcase
casez ({new_n2945_, new_n4651_})
2'b1? : new_n443_ = 1'b1;
2'b?1 : new_n443_ = 1'b1;
default : new_n443_ = 1'b0;
endcase
casez ({y[2], u[2]})
2'b00 : new_n444_ = 1'b1;
default : new_n444_ = 1'b0;
endcase
casez ({v[0], new_n82_})
2'b01 : new_n445_ = 1'b1;
default : new_n445_ = 1'b0;
endcase
casez ({new_n1174_, new_n2777_})
2'b1? : new_n446_ = 1'b1;
2'b?1 : new_n446_ = 1'b1;
default : new_n446_ = 1'b0;
endcase
casez ({new_n77_, new_n141_})
2'b01 : new_n447_ = 1'b1;
default : new_n447_ = 1'b0;
endcase
casez ({u[0], new_n152_})
2'b01 : new_n448_ = 1'b1;
default : new_n448_ = 1'b0;
endcase
casez ({new_n86_, new_n147_})
2'b11 : new_n449_ = 1'b1;
default : new_n449_ = 1'b0;
endcase
casez ({new_n97_, new_n123_})
2'b11 : new_n450_ = 1'b1;
default : new_n450_ = 1'b0;
endcase
casez ({new_n83_, new_n126_})
2'b11 : new_n451_ = 1'b1;
default : new_n451_ = 1'b0;
endcase
casez ({new_n713_, new_n265_})
2'b1? : new_n452_ = 1'b1;
2'b?1 : new_n452_ = 1'b1;
default : new_n452_ = 1'b0;
endcase
casez ({new_n1579_, new_n1099_})
2'b1? : new_n453_ = 1'b1;
2'b?1 : new_n453_ = 1'b1;
default : new_n453_ = 1'b0;
endcase
casez ({u[0], new_n163_})
2'b11 : new_n454_ = 1'b1;
default : new_n454_ = 1'b0;
endcase
casez ({y[2], new_n116_})
2'b11 : new_n455_ = 1'b1;
default : new_n455_ = 1'b0;
endcase
casez ({v[1], new_n231_})
2'b01 : new_n456_ = 1'b1;
default : new_n456_ = 1'b0;
endcase
casez ({v[2], new_n128_})
2'b01 : new_n457_ = 1'b1;
default : new_n457_ = 1'b0;
endcase
casez ({new_n81_, new_n120_})
2'b01 : new_n458_ = 1'b1;
default : new_n458_ = 1'b0;
endcase
casez ({u[2], new_n133_})
2'b01 : new_n459_ = 1'b1;
default : new_n459_ = 1'b0;
endcase
casez ({new_n77_, new_n136_})
2'b11 : new_n460_ = 1'b1;
default : new_n460_ = 1'b0;
endcase
casez ({new_n1902_, new_n268_})
2'b1? : new_n461_ = 1'b1;
2'b?1 : new_n461_ = 1'b1;
default : new_n461_ = 1'b0;
endcase
casez ({v[1], new_n106_})
2'b01 : new_n462_ = 1'b1;
default : new_n462_ = 1'b0;
endcase
casez ({new_n84_, new_n185_})
2'b11 : new_n463_ = 1'b1;
default : new_n463_ = 1'b0;
endcase
casez ({new_n80_, new_n202_})
2'b11 : new_n464_ = 1'b1;
default : new_n464_ = 1'b0;
endcase
casez ({new_n237_, new_n258_})
2'b00 : new_n465_ = 1'b1;
default : new_n465_ = 1'b0;
endcase
casez ({new_n1500_, new_n1501_})
2'b1? : new_n466_ = 1'b1;
2'b?1 : new_n466_ = 1'b1;
default : new_n466_ = 1'b0;
endcase
casez ({new_n78_, new_n361_})
2'b11 : new_n467_ = 1'b1;
default : new_n467_ = 1'b0;
endcase
casez ({new_n115_, new_n164_})
2'b11 : new_n468_ = 1'b1;
default : new_n468_ = 1'b0;
endcase
casez ({u[2], new_n98_})
2'b11 : new_n469_ = 1'b1;
default : new_n469_ = 1'b0;
endcase
casez ({new_n2684_, new_n3502_})
2'b1? : new_n470_ = 1'b1;
2'b?1 : new_n470_ = 1'b1;
default : new_n470_ = 1'b0;
endcase
casez ({new_n138_, new_n153_})
2'b11 : new_n471_ = 1'b1;
default : new_n471_ = 1'b0;
endcase
casez ({x[1], new_n357_})
2'b11 : new_n472_ = 1'b1;
default : new_n472_ = 1'b0;
endcase
casez ({v[2], new_n130_})
2'b01 : new_n473_ = 1'b1;
default : new_n473_ = 1'b0;
endcase
casez ({new_n2847_, new_n1609_})
2'b1? : new_n474_ = 1'b1;
2'b?1 : new_n474_ = 1'b1;
default : new_n474_ = 1'b0;
endcase
casez ({new_n983_, new_n3463_})
2'b1? : new_n475_ = 1'b1;
2'b?1 : new_n475_ = 1'b1;
default : new_n475_ = 1'b0;
endcase
casez ({x[2], u[0]})
2'b10 : new_n476_ = 1'b1;
default : new_n476_ = 1'b0;
endcase
casez ({new_n1632_, new_n2736_})
2'b1? : new_n477_ = 1'b1;
2'b?1 : new_n477_ = 1'b1;
default : new_n477_ = 1'b0;
endcase
casez ({new_n81_, new_n90_})
2'b01 : new_n478_ = 1'b1;
default : new_n478_ = 1'b0;
endcase
casez ({new_n955_, new_n3591_})
2'b1? : new_n479_ = 1'b1;
2'b?1 : new_n479_ = 1'b1;
default : new_n479_ = 1'b0;
endcase
casez ({y[0], new_n77_})
2'b00 : new_n480_ = 1'b1;
default : new_n480_ = 1'b0;
endcase
casez ({new_n95_, new_n141_})
2'b11 : new_n481_ = 1'b1;
default : new_n481_ = 1'b0;
endcase
casez ({new_n129_, new_n154_})
2'b11 : new_n482_ = 1'b1;
default : new_n482_ = 1'b0;
endcase
casez ({new_n86_, new_n165_})
2'b11 : new_n483_ = 1'b1;
default : new_n483_ = 1'b0;
endcase
casez ({v[1], new_n235_})
2'b01 : new_n484_ = 1'b1;
default : new_n484_ = 1'b0;
endcase
casez ({new_n269_, new_n416_})
2'b00 : new_n485_ = 1'b1;
default : new_n485_ = 1'b0;
endcase
casez ({y[0], v[2]})
2'b11 : new_n486_ = 1'b1;
default : new_n486_ = 1'b0;
endcase
casez ({y[0], v[2]})
2'b10 : new_n487_ = 1'b1;
default : new_n487_ = 1'b0;
endcase
casez ({u[2], new_n98_})
2'b01 : new_n488_ = 1'b1;
default : new_n488_ = 1'b0;
endcase
casez ({new_n80_, new_n83_})
2'b01 : new_n489_ = 1'b1;
default : new_n489_ = 1'b0;
endcase
casez ({new_n1387_, new_n2754_})
2'b1? : new_n490_ = 1'b1;
2'b?1 : new_n490_ = 1'b1;
default : new_n490_ = 1'b0;
endcase
casez ({new_n261_, new_n285_})
2'b00 : new_n491_ = 1'b1;
default : new_n491_ = 1'b0;
endcase
casez ({new_n220_, new_n247_})
2'b00 : new_n492_ = 1'b1;
default : new_n492_ = 1'b0;
endcase
casez ({y[2], new_n107_})
2'b10 : new_n493_ = 1'b1;
default : new_n493_ = 1'b0;
endcase
casez ({new_n97_, new_n116_})
2'b11 : new_n494_ = 1'b1;
default : new_n494_ = 1'b0;
endcase
casez ({v[2], new_n136_})
2'b01 : new_n495_ = 1'b1;
default : new_n495_ = 1'b0;
endcase
casez ({new_n85_, new_n146_})
2'b11 : new_n496_ = 1'b1;
default : new_n496_ = 1'b0;
endcase
casez ({x[0], new_n119_})
2'b11 : new_n497_ = 1'b1;
default : new_n497_ = 1'b0;
endcase
casez ({new_n79_, new_n138_})
2'b11 : new_n498_ = 1'b1;
default : new_n498_ = 1'b0;
endcase
casez ({new_n597_, new_n95_})
2'b1? : new_n499_ = 1'b1;
2'b?1 : new_n499_ = 1'b1;
default : new_n499_ = 1'b0;
endcase
casez ({y[1], new_n90_})
2'b11 : new_n500_ = 1'b1;
default : new_n500_ = 1'b0;
endcase
casez ({u[0], new_n163_})
2'b01 : new_n501_ = 1'b1;
default : new_n501_ = 1'b0;
endcase
casez ({new_n95_, new_n180_})
2'b11 : new_n502_ = 1'b1;
default : new_n502_ = 1'b0;
endcase
casez ({new_n79_, new_n183_})
2'b01 : new_n503_ = 1'b1;
default : new_n503_ = 1'b0;
endcase
casez ({new_n87_, new_n184_})
2'b11 : new_n504_ = 1'b1;
default : new_n504_ = 1'b0;
endcase
casez ({new_n77_, new_n130_})
2'b11 : new_n505_ = 1'b1;
default : new_n505_ = 1'b0;
endcase
casez ({new_n83_, new_n185_})
2'b11 : new_n506_ = 1'b1;
default : new_n506_ = 1'b0;
endcase
casez ({new_n1503_, new_n400_})
2'b1? : new_n507_ = 1'b1;
2'b?1 : new_n507_ = 1'b1;
default : new_n507_ = 1'b0;
endcase
casez ({x[1], new_n97_})
2'b11 : new_n508_ = 1'b1;
default : new_n508_ = 1'b0;
endcase
casez ({x[1], new_n97_})
2'b01 : new_n509_ = 1'b1;
default : new_n509_ = 1'b0;
endcase
casez ({new_n2721_, new_n145_, new_n273_})
3'b1?? : new_n510_ = 1'b1;
3'b?11 : new_n510_ = 1'b1;
default : new_n510_ = 1'b0;
endcase
casez ({new_n239_, new_n318_})
2'b00 : new_n511_ = 1'b1;
default : new_n511_ = 1'b0;
endcase
casez ({new_n3518_, new_n3513_})
2'b1? : new_n512_ = 1'b1;
2'b?1 : new_n512_ = 1'b1;
default : new_n512_ = 1'b0;
endcase
casez ({new_n148_, new_n213_, new_n1593_})
3'b11? : new_n513_ = 1'b1;
3'b??1 : new_n513_ = 1'b1;
default : new_n513_ = 1'b0;
endcase
casez ({new_n1897_, new_n3525_})
2'b1? : new_n514_ = 1'b1;
2'b?1 : new_n514_ = 1'b1;
default : new_n514_ = 1'b0;
endcase
casez ({new_n1958_, new_n92_, new_n184_})
3'b1?? : new_n515_ = 1'b1;
3'b?11 : new_n515_ = 1'b1;
default : new_n515_ = 1'b0;
endcase
casez ({new_n1339_, new_n1381_})
2'b1? : new_n516_ = 1'b1;
2'b?1 : new_n516_ = 1'b1;
default : new_n516_ = 1'b0;
endcase
casez ({u[2], new_n156_})
2'b01 : new_n517_ = 1'b1;
default : new_n517_ = 1'b0;
endcase
casez ({new_n2846_, new_n4669_})
2'b1? : new_n518_ = 1'b1;
2'b?1 : new_n518_ = 1'b1;
default : new_n518_ = 1'b0;
endcase
casez ({new_n814_, new_n3466_})
2'b1? : new_n519_ = 1'b1;
2'b?1 : new_n519_ = 1'b1;
default : new_n519_ = 1'b0;
endcase
casez ({y[2], new_n185_})
2'b11 : new_n520_ = 1'b1;
default : new_n520_ = 1'b0;
endcase
casez ({new_n118_, new_n168_})
2'b11 : new_n521_ = 1'b1;
default : new_n521_ = 1'b0;
endcase
casez ({y[0], y[1]})
2'b11 : new_n522_ = 1'b1;
default : new_n522_ = 1'b0;
endcase
casez ({new_n178_, new_n191_})
2'b00 : new_n523_ = 1'b1;
default : new_n523_ = 1'b0;
endcase
casez ({new_n94_, new_n147_})
2'b11 : new_n524_ = 1'b1;
default : new_n524_ = 1'b0;
endcase
casez ({x[0], new_n119_})
2'b01 : new_n525_ = 1'b1;
default : new_n525_ = 1'b0;
endcase
casez ({u[0], new_n124_})
2'b11 : new_n526_ = 1'b1;
default : new_n526_ = 1'b0;
endcase
casez ({new_n93_, new_n206_})
2'b11 : new_n527_ = 1'b1;
default : new_n527_ = 1'b0;
endcase
casez ({new_n157_, new_n179_})
2'b00 : new_n528_ = 1'b1;
default : new_n528_ = 1'b0;
endcase
casez ({new_n1898_, new_n457_})
2'b1? : new_n529_ = 1'b1;
2'b?1 : new_n529_ = 1'b1;
default : new_n529_ = 1'b0;
endcase
casez ({new_n94_, new_n99_})
2'b11 : new_n530_ = 1'b1;
default : new_n530_ = 1'b0;
endcase
casez ({new_n80_, new_n84_})
2'b01 : new_n531_ = 1'b1;
default : new_n531_ = 1'b0;
endcase
casez ({y[1], new_n90_})
2'b01 : new_n532_ = 1'b1;
default : new_n532_ = 1'b0;
endcase
casez ({new_n743_, new_n960_})
2'b1? : new_n533_ = 1'b1;
2'b?1 : new_n533_ = 1'b1;
default : new_n533_ = 1'b0;
endcase
casez ({new_n1940_, new_n3543_})
2'b1? : new_n534_ = 1'b1;
2'b?1 : new_n534_ = 1'b1;
default : new_n534_ = 1'b0;
endcase
casez ({new_n140_, new_n142_})
2'b11 : new_n535_ = 1'b1;
default : new_n535_ = 1'b0;
endcase
casez ({u[0], new_n143_})
2'b01 : new_n536_ = 1'b1;
default : new_n536_ = 1'b0;
endcase
casez ({new_n81_, new_n147_})
2'b11 : new_n537_ = 1'b1;
default : new_n537_ = 1'b0;
endcase
casez ({new_n89_, new_n152_})
2'b11 : new_n538_ = 1'b1;
default : new_n538_ = 1'b0;
endcase
casez ({v[1], new_n155_})
2'b11 : new_n539_ = 1'b1;
default : new_n539_ = 1'b0;
endcase
casez ({new_n115_, new_n158_})
2'b11 : new_n540_ = 1'b1;
default : new_n540_ = 1'b0;
endcase
casez ({y[2], new_n107_})
2'b00 : new_n541_ = 1'b1;
default : new_n541_ = 1'b0;
endcase
casez ({u[0], new_n124_})
2'b01 : new_n542_ = 1'b1;
default : new_n542_ = 1'b0;
endcase
casez ({new_n87_, new_n133_})
2'b11 : new_n543_ = 1'b1;
default : new_n543_ = 1'b0;
endcase
casez ({y[2], new_n185_})
2'b01 : new_n544_ = 1'b1;
default : new_n544_ = 1'b0;
endcase
casez ({new_n90_, new_n105_})
2'b11 : new_n545_ = 1'b1;
default : new_n545_ = 1'b0;
endcase
casez ({new_n83_, new_n283_})
2'b11 : new_n546_ = 1'b1;
default : new_n546_ = 1'b0;
endcase
casez ({new_n164_, new_n209_})
2'b11 : new_n547_ = 1'b1;
default : new_n547_ = 1'b0;
endcase
casez ({new_n1755_, new_n468_})
2'b1? : new_n548_ = 1'b1;
2'b?1 : new_n548_ = 1'b1;
default : new_n548_ = 1'b0;
endcase
casez ({new_n706_, v[2]})
2'b1? : new_n549_ = 1'b1;
2'b?0 : new_n549_ = 1'b1;
default : new_n549_ = 1'b0;
endcase
casez ({new_n237_, new_n347_})
2'b00 : new_n550_ = 1'b1;
default : new_n550_ = 1'b0;
endcase
casez ({x[0], new_n143_})
2'b01 : new_n551_ = 1'b1;
default : new_n551_ = 1'b0;
endcase
casez ({x[0], new_n143_})
2'b11 : new_n552_ = 1'b1;
default : new_n552_ = 1'b0;
endcase
casez ({new_n127_, new_n148_})
2'b11 : new_n553_ = 1'b1;
default : new_n553_ = 1'b0;
endcase
casez ({new_n88_, new_n152_})
2'b11 : new_n554_ = 1'b1;
default : new_n554_ = 1'b0;
endcase
casez ({new_n85_, new_n165_})
2'b11 : new_n555_ = 1'b1;
default : new_n555_ = 1'b0;
endcase
casez ({new_n87_, new_n174_})
2'b01 : new_n556_ = 1'b1;
default : new_n556_ = 1'b0;
endcase
casez ({new_n82_, new_n120_})
2'b11 : new_n557_ = 1'b1;
default : new_n557_ = 1'b0;
endcase
casez ({u[0], new_n87_})
2'b00 : new_n558_ = 1'b1;
default : new_n558_ = 1'b0;
endcase
casez ({new_n1498_, new_n4645_})
2'b1? : new_n559_ = 1'b1;
2'b?1 : new_n559_ = 1'b1;
default : new_n559_ = 1'b0;
endcase
casez ({new_n727_, new_n259_})
2'b1? : new_n560_ = 1'b1;
2'b?1 : new_n560_ = 1'b1;
default : new_n560_ = 1'b0;
endcase
casez ({new_n108_, new_n206_})
2'b11 : new_n561_ = 1'b1;
default : new_n561_ = 1'b0;
endcase
casez ({y[2], new_n277_})
2'b01 : new_n562_ = 1'b1;
default : new_n562_ = 1'b0;
endcase
casez ({new_n83_, new_n164_})
2'b11 : new_n563_ = 1'b1;
default : new_n563_ = 1'b0;
endcase
casez ({new_n86_, new_n88_})
2'b00 : new_n564_ = 1'b1;
default : new_n564_ = 1'b0;
endcase
casez ({v[1], new_n337_})
2'b01 : new_n565_ = 1'b1;
default : new_n565_ = 1'b0;
endcase
casez ({new_n1359_, new_n3462_})
2'b1? : new_n566_ = 1'b1;
2'b?1 : new_n566_ = 1'b1;
default : new_n566_ = 1'b0;
endcase
casez ({new_n1142_, new_n139_, new_n281_})
3'b1?? : new_n567_ = 1'b1;
3'b?11 : new_n567_ = 1'b1;
default : new_n567_ = 1'b0;
endcase
casez ({new_n140_, new_n198_, new_n2719_})
3'b11? : new_n568_ = 1'b1;
3'b??1 : new_n568_ = 1'b1;
default : new_n568_ = 1'b0;
endcase
casez ({new_n1021_, new_n677_})
2'b1? : new_n569_ = 1'b1;
2'b?1 : new_n569_ = 1'b1;
default : new_n569_ = 1'b0;
endcase
casez ({new_n115_, new_n266_, new_n118_, new_n342_})
4'b11?? : new_n570_ = 1'b1;
4'b??11 : new_n570_ = 1'b1;
default : new_n570_ = 1'b0;
endcase
casez ({new_n956_, u[2], new_n204_})
3'b1?? : new_n571_ = 1'b1;
3'b?01 : new_n571_ = 1'b1;
default : new_n571_ = 1'b0;
endcase
casez ({new_n1168_, new_n2763_})
2'b1? : new_n572_ = 1'b1;
2'b?1 : new_n572_ = 1'b1;
default : new_n572_ = 1'b0;
endcase
casez ({new_n115_, new_n427_, new_n118_, new_n285_})
4'b11?? : new_n573_ = 1'b1;
4'b??11 : new_n573_ = 1'b1;
default : new_n573_ = 1'b0;
endcase
casez ({new_n158_, new_n229_})
2'b00 : new_n574_ = 1'b1;
default : new_n574_ = 1'b0;
endcase
casez ({new_n131_, new_n433_, new_n213_, new_n219_})
4'b11?? : new_n575_ = 1'b1;
4'b??11 : new_n575_ = 1'b1;
default : new_n575_ = 1'b0;
endcase
casez ({new_n682_, new_n752_})
2'b1? : new_n576_ = 1'b1;
2'b?1 : new_n576_ = 1'b1;
default : new_n576_ = 1'b0;
endcase
casez ({new_n137_, new_n142_})
2'b11 : new_n577_ = 1'b1;
default : new_n577_ = 1'b0;
endcase
casez ({new_n77_, new_n147_})
2'b01 : new_n578_ = 1'b1;
default : new_n578_ = 1'b0;
endcase
casez ({new_n107_, new_n156_})
2'b01 : new_n579_ = 1'b1;
default : new_n579_ = 1'b0;
endcase
casez ({new_n137_, new_n169_})
2'b11 : new_n580_ = 1'b1;
default : new_n580_ = 1'b0;
endcase
casez ({new_n92_, new_n206_})
2'b11 : new_n581_ = 1'b1;
default : new_n581_ = 1'b0;
endcase
casez ({new_n80_, new_n238_})
2'b01 : new_n582_ = 1'b1;
default : new_n582_ = 1'b0;
endcase
casez ({y[2], new_n126_})
2'b11 : new_n583_ = 1'b1;
default : new_n583_ = 1'b0;
endcase
casez ({x[0], new_n135_})
2'b01 : new_n584_ = 1'b1;
default : new_n584_ = 1'b0;
endcase
casez ({new_n1221_, new_n2155_})
2'b1? : new_n585_ = 1'b1;
2'b?1 : new_n585_ = 1'b1;
default : new_n585_ = 1'b0;
endcase
casez ({u[2], new_n245_, new_n123_, new_n274_})
4'b01?? : new_n586_ = 1'b1;
4'b??11 : new_n586_ = 1'b1;
default : new_n586_ = 1'b0;
endcase
casez ({new_n1223_, new_n2704_})
2'b1? : new_n587_ = 1'b1;
2'b?1 : new_n587_ = 1'b1;
default : new_n587_ = 1'b0;
endcase
casez ({new_n1497_, new_n862_})
2'b1? : new_n588_ = 1'b1;
2'b?1 : new_n588_ = 1'b1;
default : new_n588_ = 1'b0;
endcase
casez ({new_n1499_, new_n2691_})
2'b1? : new_n589_ = 1'b1;
2'b?1 : new_n589_ = 1'b1;
default : new_n589_ = 1'b0;
endcase
casez ({new_n1751_, new_n3501_})
2'b1? : new_n590_ = 1'b1;
2'b?1 : new_n590_ = 1'b1;
default : new_n590_ = 1'b0;
endcase
casez ({new_n1498_, new_n1502_})
2'b1? : new_n591_ = 1'b1;
2'b?1 : new_n591_ = 1'b1;
default : new_n591_ = 1'b0;
endcase
casez ({new_n2137_, new_n1754_})
2'b1? : new_n592_ = 1'b1;
2'b?1 : new_n592_ = 1'b1;
default : new_n592_ = 1'b0;
endcase
casez ({new_n115_, new_n134_, new_n118_, new_n132_})
4'b11?? : new_n593_ = 1'b1;
4'b??11 : new_n593_ = 1'b1;
default : new_n593_ = 1'b0;
endcase
casez ({new_n1356_, new_n150_, new_n263_})
3'b1?? : new_n594_ = 1'b1;
3'b?11 : new_n594_ = 1'b1;
default : new_n594_ = 1'b0;
endcase
casez ({new_n118_, new_n263_, new_n1007_})
3'b11? : new_n595_ = 1'b1;
3'b??1 : new_n595_ = 1'b1;
default : new_n595_ = 1'b0;
endcase
casez ({new_n1748_, new_n5458_})
2'b1? : new_n596_ = 1'b1;
2'b?1 : new_n596_ = 1'b1;
default : new_n596_ = 1'b0;
endcase
casez ({y[0], v[2]})
2'b01 : new_n597_ = 1'b1;
default : new_n597_ = 1'b0;
endcase
casez ({v[0], v[2]})
2'b10 : new_n598_ = 1'b1;
default : new_n598_ = 1'b0;
endcase
casez ({v[1], new_n96_})
2'b01 : new_n599_ = 1'b1;
default : new_n599_ = 1'b0;
endcase
casez ({new_n140_, new_n169_})
2'b11 : new_n600_ = 1'b1;
default : new_n600_ = 1'b0;
endcase
casez ({new_n124_, new_n130_})
2'b11 : new_n601_ = 1'b1;
default : new_n601_ = 1'b0;
endcase
casez ({new_n89_, new_n163_})
2'b11 : new_n602_ = 1'b1;
default : new_n602_ = 1'b0;
endcase
casez ({new_n88_, new_n163_})
2'b11 : new_n603_ = 1'b1;
default : new_n603_ = 1'b0;
endcase
casez ({v[1], new_n107_})
2'b00 : new_n604_ = 1'b1;
default : new_n604_ = 1'b0;
endcase
casez ({new_n77_, new_n130_})
2'b01 : new_n605_ = 1'b1;
default : new_n605_ = 1'b0;
endcase
casez ({y[1], new_n130_})
2'b01 : new_n606_ = 1'b1;
default : new_n606_ = 1'b0;
endcase
casez ({new_n86_, new_n87_})
2'b11 : new_n607_ = 1'b1;
default : new_n607_ = 1'b0;
endcase
casez ({new_n1163_, new_n1750_})
2'b1? : new_n608_ = 1'b1;
2'b?1 : new_n608_ = 1'b1;
default : new_n608_ = 1'b0;
endcase
casez ({new_n1161_, new_n245_})
2'b1? : new_n609_ = 1'b1;
2'b?1 : new_n609_ = 1'b1;
default : new_n609_ = 1'b0;
endcase
casez ({new_n106_, new_n142_})
2'b11 : new_n610_ = 1'b1;
default : new_n610_ = 1'b0;
endcase
casez ({new_n104_, new_n271_})
2'b11 : new_n611_ = 1'b1;
default : new_n611_ = 1'b0;
endcase
casez ({new_n97_, new_n186_})
2'b11 : new_n612_ = 1'b1;
default : new_n612_ = 1'b0;
endcase
casez ({new_n84_, new_n236_})
2'b11 : new_n613_ = 1'b1;
default : new_n613_ = 1'b0;
endcase
casez ({new_n83_, new_n331_})
2'b11 : new_n614_ = 1'b1;
default : new_n614_ = 1'b0;
endcase
casez ({new_n81_, new_n437_})
2'b00 : new_n615_ = 1'b1;
default : new_n615_ = 1'b0;
endcase
casez ({x[1], new_n98_})
2'b11 : new_n616_ = 1'b1;
default : new_n616_ = 1'b0;
endcase
casez ({new_n123_, new_n154_})
2'b11 : new_n617_ = 1'b1;
default : new_n617_ = 1'b0;
endcase
casez ({y[2], new_n140_})
2'b01 : new_n618_ = 1'b1;
default : new_n618_ = 1'b0;
endcase
casez ({new_n97_, new_n107_})
2'b10 : new_n619_ = 1'b1;
default : new_n619_ = 1'b0;
endcase
casez ({new_n86_, new_n118_})
2'b11 : new_n620_ = 1'b1;
default : new_n620_ = 1'b0;
endcase
casez ({new_n1399_, new_n289_})
2'b1? : new_n621_ = 1'b1;
2'b?1 : new_n621_ = 1'b1;
default : new_n621_ = 1'b0;
endcase
casez ({new_n104_, new_n142_, new_n435_})
3'b11? : new_n622_ = 1'b1;
3'b??1 : new_n622_ = 1'b1;
default : new_n622_ = 1'b0;
endcase
casez ({v[1], new_n157_})
2'b11 : new_n623_ = 1'b1;
default : new_n623_ = 1'b0;
endcase
casez ({new_n83_, new_n236_})
2'b11 : new_n624_ = 1'b1;
default : new_n624_ = 1'b0;
endcase
casez ({new_n93_, new_n245_})
2'b11 : new_n625_ = 1'b1;
default : new_n625_ = 1'b0;
endcase
casez ({new_n117_, new_n142_})
2'b11 : new_n626_ = 1'b1;
default : new_n626_ = 1'b0;
endcase
casez ({new_n2764_, u[2], new_n187_})
3'b1?? : new_n627_ = 1'b1;
3'b?01 : new_n627_ = 1'b1;
default : new_n627_ = 1'b0;
endcase
casez ({new_n167_, new_n208_})
2'b00 : new_n628_ = 1'b1;
default : new_n628_ = 1'b0;
endcase
casez ({new_n123_, new_n213_})
2'b00 : new_n629_ = 1'b1;
default : new_n629_ = 1'b0;
endcase
casez ({new_n176_, new_n258_})
2'b00 : new_n630_ = 1'b1;
default : new_n630_ = 1'b0;
endcase
casez ({new_n124_, new_n165_})
2'b11 : new_n631_ = 1'b1;
default : new_n631_ = 1'b0;
endcase
casez ({new_n96_, new_n228_})
2'b11 : new_n632_ = 1'b1;
default : new_n632_ = 1'b0;
endcase
casez ({v[2], new_n130_})
2'b11 : new_n633_ = 1'b1;
default : new_n633_ = 1'b0;
endcase
casez ({new_n94_, new_n165_})
2'b11 : new_n634_ = 1'b1;
default : new_n634_ = 1'b0;
endcase
casez ({new_n109_, new_n170_})
2'b01 : new_n635_ = 1'b1;
default : new_n635_ = 1'b0;
endcase
casez ({y[2], new_n129_})
2'b01 : new_n636_ = 1'b1;
default : new_n636_ = 1'b0;
endcase
casez ({new_n97_, new_n129_})
2'b11 : new_n637_ = 1'b1;
default : new_n637_ = 1'b0;
endcase
casez ({new_n86_, new_n131_})
2'b11 : new_n638_ = 1'b1;
default : new_n638_ = 1'b0;
endcase
casez ({new_n86_, new_n139_})
2'b11 : new_n639_ = 1'b1;
default : new_n639_ = 1'b0;
endcase
casez ({new_n137_, new_n148_, new_n535_})
3'b11? : new_n640_ = 1'b1;
3'b??1 : new_n640_ = 1'b1;
default : new_n640_ = 1'b0;
endcase
casez ({new_n202_, new_n539_})
2'b00 : new_n641_ = 1'b1;
default : new_n641_ = 1'b0;
endcase
casez ({new_n112_, new_n142_})
2'b11 : new_n642_ = 1'b1;
default : new_n642_ = 1'b0;
endcase
casez ({new_n110_, new_n142_})
2'b11 : new_n643_ = 1'b1;
default : new_n643_ = 1'b0;
endcase
casez ({new_n83_, new_n286_})
2'b11 : new_n644_ = 1'b1;
default : new_n644_ = 1'b0;
endcase
casez ({new_n84_, new_n292_})
2'b11 : new_n645_ = 1'b1;
default : new_n645_ = 1'b0;
endcase
casez ({x[0], new_n310_})
2'b11 : new_n646_ = 1'b1;
default : new_n646_ = 1'b0;
endcase
casez ({new_n115_, new_n179_})
2'b11 : new_n647_ = 1'b1;
default : new_n647_ = 1'b0;
endcase
casez ({y[0], new_n105_})
2'b11 : new_n648_ = 1'b1;
default : new_n648_ = 1'b0;
endcase
casez ({y[0], new_n421_})
2'b01 : new_n649_ = 1'b1;
default : new_n649_ = 1'b0;
endcase
casez ({new_n426_, new_n496_})
2'b00 : new_n650_ = 1'b1;
default : new_n650_ = 1'b0;
endcase
casez ({new_n92_, new_n280_, new_n131_, new_n246_})
4'b11?? : new_n651_ = 1'b1;
4'b??11 : new_n651_ = 1'b1;
default : new_n651_ = 1'b0;
endcase
casez ({new_n83_, new_n168_, new_n84_, new_n164_})
4'b11?? : new_n652_ = 1'b1;
4'b??11 : new_n652_ = 1'b1;
default : new_n652_ = 1'b0;
endcase
casez ({x[0], new_n168_})
2'b01 : new_n653_ = 1'b1;
default : new_n653_ = 1'b0;
endcase
casez ({new_n82_, new_n98_})
2'b01 : new_n654_ = 1'b1;
default : new_n654_ = 1'b0;
endcase
casez ({new_n2683_, new_n129_, new_n142_})
3'b1?? : new_n655_ = 1'b1;
3'b?11 : new_n655_ = 1'b1;
default : new_n655_ = 1'b0;
endcase
casez ({new_n89_, new_n103_, new_n160_})
3'b10? : new_n656_ = 1'b1;
3'b??1 : new_n656_ = 1'b1;
default : new_n656_ = 1'b0;
endcase
casez ({new_n3484_, new_n2686_})
2'b1? : new_n657_ = 1'b1;
2'b?1 : new_n657_ = 1'b1;
default : new_n657_ = 1'b0;
endcase
casez ({new_n118_, new_n307_, new_n162_, new_n266_})
4'b11?? : new_n658_ = 1'b1;
4'b??11 : new_n658_ = 1'b1;
default : new_n658_ = 1'b0;
endcase
casez ({new_n95_, new_n222_})
2'b00 : new_n659_ = 1'b1;
default : new_n659_ = 1'b0;
endcase
casez ({new_n1350_, new_n154_, new_n160_})
3'b1?? : new_n660_ = 1'b1;
3'b?11 : new_n660_ = 1'b1;
default : new_n660_ = 1'b0;
endcase
casez ({new_n144_, new_n317_, new_n3499_})
3'b11? : new_n661_ = 1'b1;
3'b??1 : new_n661_ = 1'b1;
default : new_n661_ = 1'b0;
endcase
casez ({new_n3595_, new_n1904_})
2'b1? : new_n662_ = 1'b1;
2'b?1 : new_n662_ = 1'b1;
default : new_n662_ = 1'b0;
endcase
casez ({new_n2698_, new_n2727_})
2'b1? : new_n663_ = 1'b1;
2'b?1 : new_n663_ = 1'b1;
default : new_n663_ = 1'b0;
endcase
casez ({new_n1368_, new_n1117_})
2'b1? : new_n664_ = 1'b1;
2'b?1 : new_n664_ = 1'b1;
default : new_n664_ = 1'b0;
endcase
casez ({new_n1354_, new_n2735_})
2'b1? : new_n665_ = 1'b1;
2'b?1 : new_n665_ = 1'b1;
default : new_n665_ = 1'b0;
endcase
casez ({new_n153_, new_n210_, new_n3528_})
3'b11? : new_n666_ = 1'b1;
3'b??1 : new_n666_ = 1'b1;
default : new_n666_ = 1'b0;
endcase
casez ({new_n3531_, new_n1011_})
2'b1? : new_n667_ = 1'b1;
2'b?1 : new_n667_ = 1'b1;
default : new_n667_ = 1'b0;
endcase
casez ({new_n127_, new_n154_})
2'b11 : new_n668_ = 1'b1;
default : new_n668_ = 1'b0;
endcase
casez ({x[1], new_n156_})
2'b11 : new_n669_ = 1'b1;
default : new_n669_ = 1'b0;
endcase
casez ({new_n4652_, new_n1342_})
2'b1? : new_n670_ = 1'b1;
2'b?1 : new_n670_ = 1'b1;
default : new_n670_ = 1'b0;
endcase
casez ({new_n109_, new_n156_})
2'b01 : new_n671_ = 1'b1;
default : new_n671_ = 1'b0;
endcase
casez ({v[2], new_n120_})
2'b11 : new_n672_ = 1'b1;
default : new_n672_ = 1'b0;
endcase
casez ({v[1], new_n145_})
2'b11 : new_n673_ = 1'b1;
default : new_n673_ = 1'b0;
endcase
casez ({x[0], new_n152_})
2'b01 : new_n674_ = 1'b1;
default : new_n674_ = 1'b0;
endcase
casez ({u[2], new_n159_})
2'b01 : new_n675_ = 1'b1;
default : new_n675_ = 1'b0;
endcase
casez ({new_n80_, new_n182_})
2'b01 : new_n676_ = 1'b1;
default : new_n676_ = 1'b0;
endcase
casez ({new_n131_, new_n201_})
2'b11 : new_n677_ = 1'b1;
default : new_n677_ = 1'b0;
endcase
casez ({new_n127_, new_n191_})
2'b11 : new_n678_ = 1'b1;
default : new_n678_ = 1'b0;
endcase
casez ({new_n88_, new_n119_})
2'b11 : new_n679_ = 1'b1;
default : new_n679_ = 1'b0;
endcase
casez ({new_n88_, new_n124_})
2'b11 : new_n680_ = 1'b1;
default : new_n680_ = 1'b0;
endcase
casez ({new_n101_, new_n124_})
2'b11 : new_n681_ = 1'b1;
default : new_n681_ = 1'b0;
endcase
casez ({u[0], new_n135_})
2'b01 : new_n682_ = 1'b1;
default : new_n682_ = 1'b0;
endcase
casez ({y[2], new_n137_})
2'b11 : new_n683_ = 1'b1;
default : new_n683_ = 1'b0;
endcase
casez ({new_n4644_, new_n3556_})
2'b1? : new_n684_ = 1'b1;
2'b?1 : new_n684_ = 1'b1;
default : new_n684_ = 1'b0;
endcase
casez ({v[1], new_n286_, new_n1144_})
3'b01? : new_n685_ = 1'b1;
3'b??1 : new_n685_ = 1'b1;
default : new_n685_ = 1'b0;
endcase
casez ({new_n1400_, new_n539_})
2'b1? : new_n686_ = 1'b1;
2'b?1 : new_n686_ = 1'b1;
default : new_n686_ = 1'b0;
endcase
casez ({new_n983_, new_n3562_})
2'b1? : new_n687_ = 1'b1;
2'b?1 : new_n687_ = 1'b1;
default : new_n687_ = 1'b0;
endcase
casez ({y[2], new_n336_, new_n1587_})
3'b11? : new_n688_ = 1'b1;
3'b??1 : new_n688_ = 1'b1;
default : new_n688_ = 1'b0;
endcase
casez ({y[2], new_n350_, new_n153_, new_n174_})
4'b11?? : new_n689_ = 1'b1;
4'b??11 : new_n689_ = 1'b1;
default : new_n689_ = 1'b0;
endcase
casez ({new_n1478_, new_n1015_})
2'b1? : new_n690_ = 1'b1;
2'b?1 : new_n690_ = 1'b1;
default : new_n690_ = 1'b0;
endcase
casez ({new_n985_, new_n2728_})
2'b1? : new_n691_ = 1'b1;
2'b?1 : new_n691_ = 1'b1;
default : new_n691_ = 1'b0;
endcase
casez ({new_n2147_, new_n3468_})
2'b1? : new_n692_ = 1'b1;
2'b?1 : new_n692_ = 1'b1;
default : new_n692_ = 1'b0;
endcase
casez ({new_n2840_, new_n82_, new_n199_})
3'b1?? : new_n693_ = 1'b1;
3'b?11 : new_n693_ = 1'b1;
default : new_n693_ = 1'b0;
endcase
casez ({new_n447_, new_n460_})
2'b00 : new_n694_ = 1'b1;
default : new_n694_ = 1'b0;
endcase
casez ({new_n84_, new_n171_})
2'b11 : new_n695_ = 1'b1;
default : new_n695_ = 1'b0;
endcase
casez ({new_n118_, new_n175_})
2'b11 : new_n696_ = 1'b1;
default : new_n696_ = 1'b0;
endcase
casez ({new_n84_, new_n175_})
2'b11 : new_n697_ = 1'b1;
default : new_n697_ = 1'b0;
endcase
casez ({new_n97_, new_n185_})
2'b11 : new_n698_ = 1'b1;
default : new_n698_ = 1'b0;
endcase
casez ({new_n111_, new_n206_})
2'b11 : new_n699_ = 1'b1;
default : new_n699_ = 1'b0;
endcase
casez ({new_n80_, new_n188_, new_n139_, new_n155_})
4'b11?? : new_n700_ = 1'b1;
4'b??11 : new_n700_ = 1'b1;
default : new_n700_ = 1'b0;
endcase
casez ({new_n984_, new_n355_})
2'b1? : new_n701_ = 1'b1;
2'b?1 : new_n701_ = 1'b1;
default : new_n701_ = 1'b0;
endcase
casez ({new_n115_, new_n239_, new_n470_})
3'b11? : new_n702_ = 1'b1;
3'b??1 : new_n702_ = 1'b1;
default : new_n702_ = 1'b0;
endcase
casez ({new_n84_, new_n168_})
2'b11 : new_n703_ = 1'b1;
default : new_n703_ = 1'b0;
endcase
casez ({new_n83_, new_n246_})
2'b11 : new_n704_ = 1'b1;
default : new_n704_ = 1'b0;
endcase
casez ({new_n4605_, new_n519_})
2'b1? : new_n705_ = 1'b1;
2'b?1 : new_n705_ = 1'b1;
default : new_n705_ = 1'b0;
endcase
casez ({y[0], y[1]})
2'b00 : new_n706_ = 1'b1;
default : new_n706_ = 1'b0;
endcase
casez ({new_n217_, new_n307_})
2'b00 : new_n707_ = 1'b1;
default : new_n707_ = 1'b0;
endcase
casez ({new_n1023_, new_n182_})
2'b1? : new_n708_ = 1'b1;
2'b?1 : new_n708_ = 1'b1;
default : new_n708_ = 1'b0;
endcase
casez ({new_n251_, new_n293_})
2'b00 : new_n709_ = 1'b1;
default : new_n709_ = 1'b0;
endcase
casez ({new_n137_, new_n260_})
2'b11 : new_n710_ = 1'b1;
default : new_n710_ = 1'b0;
endcase
casez ({new_n124_, new_n147_})
2'b11 : new_n711_ = 1'b1;
default : new_n711_ = 1'b0;
endcase
casez ({y[2], new_n109_})
2'b00 : new_n712_ = 1'b1;
default : new_n712_ = 1'b0;
endcase
casez ({x[0], new_n152_})
2'b11 : new_n713_ = 1'b1;
default : new_n713_ = 1'b0;
endcase
casez ({x[1], new_n161_})
2'b01 : new_n714_ = 1'b1;
default : new_n714_ = 1'b0;
endcase
casez ({v[1], new_n173_})
2'b11 : new_n715_ = 1'b1;
default : new_n715_ = 1'b0;
endcase
casez ({new_n89_, new_n119_})
2'b11 : new_n716_ = 1'b1;
default : new_n716_ = 1'b0;
endcase
casez ({y[2], new_n129_})
2'b11 : new_n717_ = 1'b1;
default : new_n717_ = 1'b0;
endcase
casez ({new_n103_, new_n131_})
2'b11 : new_n718_ = 1'b1;
default : new_n718_ = 1'b0;
endcase
casez ({new_n98_, new_n109_})
2'b10 : new_n719_ = 1'b1;
default : new_n719_ = 1'b0;
endcase
casez ({new_n185_, new_n498_})
2'b00 : new_n720_ = 1'b1;
default : new_n720_ = 1'b0;
endcase
casez ({new_n292_, new_n472_})
2'b00 : new_n721_ = 1'b1;
default : new_n721_ = 1'b0;
endcase
casez ({new_n84_, new_n157_})
2'b11 : new_n722_ = 1'b1;
default : new_n722_ = 1'b0;
endcase
casez ({new_n103_, new_n290_})
2'b11 : new_n723_ = 1'b1;
default : new_n723_ = 1'b0;
endcase
casez ({x[0], new_n294_})
2'b01 : new_n724_ = 1'b1;
default : new_n724_ = 1'b0;
endcase
casez ({new_n81_, new_n308_})
2'b11 : new_n725_ = 1'b1;
default : new_n725_ = 1'b0;
endcase
casez ({x[0], new_n345_})
2'b11 : new_n726_ = 1'b1;
default : new_n726_ = 1'b0;
endcase
casez ({new_n83_, new_n157_})
2'b11 : new_n727_ = 1'b1;
default : new_n727_ = 1'b0;
endcase
casez ({x[1], y[2]})
2'b11 : new_n728_ = 1'b1;
default : new_n728_ = 1'b0;
endcase
casez ({u[2], new_n234_})
2'b01 : new_n729_ = 1'b1;
default : new_n729_ = 1'b0;
endcase
casez ({u[0], new_n103_})
2'b01 : new_n730_ = 1'b1;
default : new_n730_ = 1'b0;
endcase
casez ({new_n2870_, new_n4663_})
2'b1? : new_n731_ = 1'b1;
2'b?1 : new_n731_ = 1'b1;
default : new_n731_ = 1'b0;
endcase
casez ({new_n3493_, new_n2685_})
2'b1? : new_n732_ = 1'b1;
2'b?1 : new_n732_ = 1'b1;
default : new_n732_ = 1'b0;
endcase
casez ({new_n3552_, new_n565_})
2'b1? : new_n733_ = 1'b1;
2'b?1 : new_n733_ = 1'b1;
default : new_n733_ = 1'b0;
endcase
casez ({new_n79_, new_n166_})
2'b01 : new_n734_ = 1'b1;
default : new_n734_ = 1'b0;
endcase
casez ({new_n127_, new_n182_})
2'b11 : new_n735_ = 1'b1;
default : new_n735_ = 1'b0;
endcase
casez ({new_n245_, new_n497_, new_n250_, new_n735_})
4'b11?? : new_n736_ = 1'b1;
4'b??11 : new_n736_ = 1'b1;
default : new_n736_ = 1'b0;
endcase
casez ({new_n191_, new_n198_})
2'b11 : new_n737_ = 1'b1;
default : new_n737_ = 1'b0;
endcase
casez ({new_n129_, new_n212_})
2'b11 : new_n738_ = 1'b1;
default : new_n738_ = 1'b0;
endcase
casez ({new_n93_, new_n208_})
2'b01 : new_n739_ = 1'b1;
default : new_n739_ = 1'b0;
endcase
casez ({new_n115_, new_n230_})
2'b11 : new_n740_ = 1'b1;
default : new_n740_ = 1'b0;
endcase
casez ({new_n104_, new_n141_})
2'b11 : new_n741_ = 1'b1;
default : new_n741_ = 1'b0;
endcase
casez ({new_n98_, new_n143_})
2'b11 : new_n742_ = 1'b1;
default : new_n742_ = 1'b0;
endcase
casez ({v[1], new_n144_})
2'b11 : new_n743_ = 1'b1;
default : new_n743_ = 1'b0;
endcase
casez ({new_n95_, new_n147_})
2'b11 : new_n744_ = 1'b1;
default : new_n744_ = 1'b0;
endcase
casez ({new_n89_, new_n156_})
2'b11 : new_n745_ = 1'b1;
default : new_n745_ = 1'b0;
endcase
casez ({new_n123_, new_n158_})
2'b11 : new_n746_ = 1'b1;
default : new_n746_ = 1'b0;
endcase
casez ({u[2], new_n161_})
2'b01 : new_n747_ = 1'b1;
default : new_n747_ = 1'b0;
endcase
casez ({new_n95_, new_n165_})
2'b11 : new_n748_ = 1'b1;
default : new_n748_ = 1'b0;
endcase
casez ({v[1], new_n126_})
2'b01 : new_n749_ = 1'b1;
default : new_n749_ = 1'b0;
endcase
casez ({new_n80_, new_n128_})
2'b11 : new_n750_ = 1'b1;
default : new_n750_ = 1'b0;
endcase
casez ({u[0], new_n116_})
2'b01 : new_n751_ = 1'b1;
default : new_n751_ = 1'b0;
endcase
casez ({new_n85_, new_n87_})
2'b10 : new_n752_ = 1'b1;
default : new_n752_ = 1'b0;
endcase
casez ({new_n202_, new_n311_})
2'b00 : new_n753_ = 1'b1;
default : new_n753_ = 1'b0;
endcase
casez ({new_n79_, new_n253_})
2'b11 : new_n754_ = 1'b1;
default : new_n754_ = 1'b0;
endcase
casez ({x[0], new_n295_})
2'b01 : new_n755_ = 1'b1;
default : new_n755_ = 1'b0;
endcase
casez ({v[1], new_n185_})
2'b01 : new_n756_ = 1'b1;
default : new_n756_ = 1'b0;
endcase
casez ({new_n102_, new_n130_})
2'b11 : new_n757_ = 1'b1;
default : new_n757_ = 1'b0;
endcase
casez ({new_n367_, new_n506_})
2'b00 : new_n758_ = 1'b1;
default : new_n758_ = 1'b0;
endcase
casez ({new_n471_, new_n520_})
2'b00 : new_n759_ = 1'b1;
default : new_n759_ = 1'b0;
endcase
casez ({new_n139_, new_n164_})
2'b11 : new_n760_ = 1'b1;
default : new_n760_ = 1'b0;
endcase
casez ({new_n468_, new_n521_})
2'b00 : new_n761_ = 1'b1;
default : new_n761_ = 1'b0;
endcase
casez ({new_n125_, new_n206_})
2'b11 : new_n762_ = 1'b1;
default : new_n762_ = 1'b0;
endcase
casez ({new_n2950_, new_n89_})
2'b1? : new_n763_ = 1'b1;
2'b?1 : new_n763_ = 1'b1;
default : new_n763_ = 1'b0;
endcase
casez ({y[0], new_n82_})
2'b10 : new_n764_ = 1'b1;
default : new_n764_ = 1'b0;
endcase
casez ({new_n85_, new_n96_})
2'b01 : new_n765_ = 1'b1;
default : new_n765_ = 1'b0;
endcase
casez ({new_n96_, new_n104_})
2'b11 : new_n766_ = 1'b1;
default : new_n766_ = 1'b0;
endcase
casez ({new_n234_, new_n411_})
2'b11 : new_n767_ = 1'b1;
default : new_n767_ = 1'b0;
endcase
casez ({new_n82_, new_n89_})
2'b11 : new_n768_ = 1'b1;
default : new_n768_ = 1'b0;
endcase
casez ({new_n1646_, new_n2756_})
2'b1? : new_n769_ = 1'b1;
2'b?1 : new_n769_ = 1'b1;
default : new_n769_ = 1'b0;
endcase
casez ({new_n1395_, new_n116_})
2'b1? : new_n770_ = 1'b1;
2'b?1 : new_n770_ = 1'b1;
default : new_n770_ = 1'b0;
endcase
casez ({new_n2771_, v[1], new_n213_})
3'b1?? : new_n771_ = 1'b1;
3'b?11 : new_n771_ = 1'b1;
default : new_n771_ = 1'b0;
endcase
casez ({y[2], new_n306_, new_n386_})
3'b11? : new_n772_ = 1'b1;
3'b0?1 : new_n772_ = 1'b1;
default : new_n772_ = 1'b0;
endcase
casez ({new_n2753_, new_n1146_})
2'b1? : new_n773_ = 1'b1;
2'b?1 : new_n773_ = 1'b1;
default : new_n773_ = 1'b0;
endcase
casez ({new_n170_, new_n224_})
2'b00 : new_n774_ = 1'b1;
default : new_n774_ = 1'b0;
endcase
casez ({new_n231_, new_n260_})
2'b11 : new_n775_ = 1'b1;
default : new_n775_ = 1'b0;
endcase
casez ({new_n77_, new_n147_})
2'b11 : new_n776_ = 1'b1;
default : new_n776_ = 1'b0;
endcase
casez ({new_n138_, new_n154_})
2'b11 : new_n777_ = 1'b1;
default : new_n777_ = 1'b0;
endcase
casez ({new_n129_, new_n287_})
2'b11 : new_n778_ = 1'b1;
default : new_n778_ = 1'b0;
endcase
casez ({new_n118_, new_n170_})
2'b11 : new_n779_ = 1'b1;
default : new_n779_ = 1'b0;
endcase
casez ({new_n148_, new_n205_})
2'b11 : new_n780_ = 1'b1;
default : new_n780_ = 1'b0;
endcase
casez ({u[2], new_n206_})
2'b01 : new_n781_ = 1'b1;
default : new_n781_ = 1'b0;
endcase
casez ({new_n123_, new_n219_})
2'b11 : new_n782_ = 1'b1;
default : new_n782_ = 1'b0;
endcase
casez ({y[2], new_n109_})
2'b10 : new_n783_ = 1'b1;
default : new_n783_ = 1'b0;
endcase
casez ({new_n169_, new_n231_})
2'b11 : new_n784_ = 1'b1;
default : new_n784_ = 1'b0;
endcase
casez ({new_n182_, new_n243_})
2'b11 : new_n785_ = 1'b1;
default : new_n785_ = 1'b0;
endcase
casez ({new_n77_, new_n136_})
2'b01 : new_n786_ = 1'b1;
default : new_n786_ = 1'b0;
endcase
casez ({new_n97_, new_n247_})
2'b11 : new_n787_ = 1'b1;
default : new_n787_ = 1'b0;
endcase
casez ({new_n138_, new_n142_})
2'b11 : new_n788_ = 1'b1;
default : new_n788_ = 1'b0;
endcase
casez ({new_n94_, new_n148_})
2'b11 : new_n789_ = 1'b1;
default : new_n789_ = 1'b0;
endcase
casez ({new_n103_, new_n154_})
2'b11 : new_n790_ = 1'b1;
default : new_n790_ = 1'b0;
endcase
casez ({new_n81_, new_n180_})
2'b11 : new_n791_ = 1'b1;
default : new_n791_ = 1'b0;
endcase
casez ({y[2], new_n189_})
2'b01 : new_n792_ = 1'b1;
default : new_n792_ = 1'b0;
endcase
casez ({u[2], new_n191_})
2'b01 : new_n793_ = 1'b1;
default : new_n793_ = 1'b0;
endcase
casez ({new_n79_, new_n199_})
2'b01 : new_n794_ = 1'b1;
default : new_n794_ = 1'b0;
endcase
casez ({u[2], new_n208_})
2'b11 : new_n795_ = 1'b1;
default : new_n795_ = 1'b0;
endcase
casez ({new_n98_, new_n107_})
2'b10 : new_n796_ = 1'b1;
default : new_n796_ = 1'b0;
endcase
casez ({new_n80_, new_n223_})
2'b01 : new_n797_ = 1'b1;
default : new_n797_ = 1'b0;
endcase
casez ({new_n85_, new_n131_})
2'b11 : new_n798_ = 1'b1;
default : new_n798_ = 1'b0;
endcase
casez ({x[0], new_n133_})
2'b11 : new_n799_ = 1'b1;
default : new_n799_ = 1'b0;
endcase
casez ({y[2], new_n137_})
2'b01 : new_n800_ = 1'b1;
default : new_n800_ = 1'b0;
endcase
casez ({new_n265_, new_n525_})
2'b00 : new_n801_ = 1'b1;
default : new_n801_ = 1'b0;
endcase
casez ({new_n1720_, new_n543_})
2'b1? : new_n802_ = 1'b1;
2'b?1 : new_n802_ = 1'b1;
default : new_n802_ = 1'b0;
endcase
casez ({new_n2715_, new_n335_})
2'b1? : new_n803_ = 1'b1;
2'b?1 : new_n803_ = 1'b1;
default : new_n803_ = 1'b0;
endcase
casez ({new_n1461_, new_n639_})
2'b1? : new_n804_ = 1'b1;
2'b?1 : new_n804_ = 1'b1;
default : new_n804_ = 1'b0;
endcase
casez ({new_n236_, new_n350_})
2'b00 : new_n805_ = 1'b1;
default : new_n805_ = 1'b0;
endcase
casez ({new_n81_, new_n251_, new_n4668_})
3'b11? : new_n806_ = 1'b1;
3'b??1 : new_n806_ = 1'b1;
default : new_n806_ = 1'b0;
endcase
casez ({new_n83_, new_n121_})
2'b11 : new_n807_ = 1'b1;
default : new_n807_ = 1'b0;
endcase
casez ({new_n80_, new_n253_})
2'b11 : new_n808_ = 1'b1;
default : new_n808_ = 1'b0;
endcase
casez ({new_n104_, new_n290_})
2'b11 : new_n809_ = 1'b1;
default : new_n809_ = 1'b0;
endcase
casez ({new_n83_, new_n171_})
2'b11 : new_n810_ = 1'b1;
default : new_n810_ = 1'b0;
endcase
casez ({new_n80_, new_n303_})
2'b11 : new_n811_ = 1'b1;
default : new_n811_ = 1'b0;
endcase
casez ({new_n83_, new_n175_})
2'b11 : new_n812_ = 1'b1;
default : new_n812_ = 1'b0;
endcase
casez ({new_n103_, new_n339_})
2'b11 : new_n813_ = 1'b1;
default : new_n813_ = 1'b0;
endcase
casez ({new_n79_, new_n202_})
2'b11 : new_n814_ = 1'b1;
default : new_n814_ = 1'b0;
endcase
casez ({new_n83_, new_n225_})
2'b11 : new_n815_ = 1'b1;
default : new_n815_ = 1'b0;
endcase
casez ({new_n115_, new_n121_})
2'b11 : new_n816_ = 1'b1;
default : new_n816_ = 1'b0;
endcase
casez ({new_n1138_, new_n644_})
2'b1? : new_n817_ = 1'b1;
2'b?1 : new_n817_ = 1'b1;
default : new_n817_ = 1'b0;
endcase
casez ({new_n79_, new_n409_, new_n5458_})
3'b10? : new_n818_ = 1'b1;
3'b??1 : new_n818_ = 1'b1;
default : new_n818_ = 1'b0;
endcase
casez ({new_n79_, new_n270_})
2'b11 : new_n819_ = 1'b1;
default : new_n819_ = 1'b0;
endcase
casez ({new_n4657_, new_n559_})
2'b1? : new_n820_ = 1'b1;
2'b?1 : new_n820_ = 1'b1;
default : new_n820_ = 1'b0;
endcase
casez ({new_n94_, new_n97_})
2'b11 : new_n821_ = 1'b1;
default : new_n821_ = 1'b0;
endcase
casez ({y[0], new_n81_})
2'b00 : new_n822_ = 1'b1;
default : new_n822_ = 1'b0;
endcase
casez ({new_n3479_, new_n1636_})
2'b1? : new_n823_ = 1'b1;
2'b?1 : new_n823_ = 1'b1;
default : new_n823_ = 1'b0;
endcase
casez ({new_n1607_, new_n1361_})
2'b1? : new_n824_ = 1'b1;
2'b?1 : new_n824_ = 1'b1;
default : new_n824_ = 1'b0;
endcase
casez ({new_n2772_, new_n153_, new_n500_})
3'b1?? : new_n825_ = 1'b1;
3'b?11 : new_n825_ = 1'b1;
default : new_n825_ = 1'b0;
endcase
casez ({new_n115_, new_n486_, new_n118_, new_n262_})
4'b11?? : new_n826_ = 1'b1;
4'b??11 : new_n826_ = 1'b1;
default : new_n826_ = 1'b0;
endcase
casez ({new_n167_, new_n264_, new_n1918_})
3'b11? : new_n827_ = 1'b1;
3'b??1 : new_n827_ = 1'b1;
default : new_n827_ = 1'b0;
endcase
casez ({new_n144_, new_n162_, new_n148_, new_n532_})
4'b11?? : new_n828_ = 1'b1;
4'b??11 : new_n828_ = 1'b1;
default : new_n828_ = 1'b0;
endcase
casez ({new_n2504_, new_n285_})
2'b1? : new_n829_ = 1'b1;
2'b?1 : new_n829_ = 1'b1;
default : new_n829_ = 1'b0;
endcase
casez ({new_n118_, new_n155_, new_n2709_})
3'b11? : new_n830_ = 1'b1;
3'b??1 : new_n830_ = 1'b1;
default : new_n830_ = 1'b0;
endcase
casez ({new_n241_, new_n313_, new_n249_, new_n261_})
4'b11?? : new_n831_ = 1'b1;
4'b??11 : new_n831_ = 1'b1;
default : new_n831_ = 1'b0;
endcase
casez ({new_n3370_, new_n279_, new_n316_})
3'b1?? : new_n832_ = 1'b1;
3'b?11 : new_n832_ = 1'b1;
default : new_n832_ = 1'b0;
endcase
casez ({new_n155_, new_n321_, new_n213_, new_n317_})
4'b11?? : new_n833_ = 1'b1;
4'b??11 : new_n833_ = 1'b1;
default : new_n833_ = 1'b0;
endcase
casez ({new_n153_, new_n201_, new_n182_, new_n328_})
4'b11?? : new_n834_ = 1'b1;
4'b??11 : new_n834_ = 1'b1;
default : new_n834_ = 1'b0;
endcase
casez ({new_n1178_, new_n3401_})
2'b1? : new_n835_ = 1'b1;
2'b?1 : new_n835_ = 1'b1;
default : new_n835_ = 1'b0;
endcase
casez ({new_n2587_, new_n173_, new_n363_})
3'b1?? : new_n836_ = 1'b1;
3'b?11 : new_n836_ = 1'b1;
default : new_n836_ = 1'b0;
endcase
casez ({new_n1140_, new_n150_, new_n205_})
3'b1?? : new_n837_ = 1'b1;
3'b?11 : new_n837_ = 1'b1;
default : new_n837_ = 1'b0;
endcase
casez ({new_n1914_, new_n1912_})
2'b1? : new_n838_ = 1'b1;
2'b?1 : new_n838_ = 1'b1;
default : new_n838_ = 1'b0;
endcase
casez ({new_n3595_, new_n2731_})
2'b1? : new_n839_ = 1'b1;
2'b?1 : new_n839_ = 1'b1;
default : new_n839_ = 1'b0;
endcase
casez ({new_n2690_, new_n2737_})
2'b1? : new_n840_ = 1'b1;
2'b?1 : new_n840_ = 1'b1;
default : new_n840_ = 1'b0;
endcase
casez ({new_n115_, new_n140_, new_n153_, new_n218_})
4'b11?? : new_n841_ = 1'b1;
4'b??11 : new_n841_ = 1'b1;
default : new_n841_ = 1'b0;
endcase
casez ({new_n1925_, new_n1102_})
2'b1? : new_n842_ = 1'b1;
2'b?1 : new_n842_ = 1'b1;
default : new_n842_ = 1'b0;
endcase
casez ({new_n1372_, new_n139_, new_n226_})
3'b1?? : new_n843_ = 1'b1;
3'b?11 : new_n843_ = 1'b1;
default : new_n843_ = 1'b0;
endcase
casez ({new_n139_, new_n427_, new_n3356_})
3'b11? : new_n844_ = 1'b1;
3'b??1 : new_n844_ = 1'b1;
default : new_n844_ = 1'b0;
endcase
casez ({new_n3464_, new_n92_, new_n230_})
3'b1?? : new_n845_ = 1'b1;
3'b?11 : new_n845_ = 1'b1;
default : new_n845_ = 1'b0;
endcase
casez ({new_n3551_, new_n3563_})
2'b1? : new_n846_ = 1'b1;
2'b?1 : new_n846_ = 1'b1;
default : new_n846_ = 1'b0;
endcase
casez ({new_n150_, new_n438_, new_n190_, new_n207_})
4'b11?? : new_n847_ = 1'b1;
4'b??11 : new_n847_ = 1'b1;
default : new_n847_ = 1'b0;
endcase
casez ({new_n115_, new_n137_, new_n153_, new_n226_})
4'b11?? : new_n848_ = 1'b1;
4'b??11 : new_n848_ = 1'b1;
default : new_n848_ = 1'b0;
endcase
casez ({new_n139_, new_n240_, new_n3425_})
3'b11? : new_n849_ = 1'b1;
3'b??1 : new_n849_ = 1'b1;
default : new_n849_ = 1'b0;
endcase
casez ({new_n131_, new_n239_, new_n189_, new_n241_})
4'b11?? : new_n850_ = 1'b1;
4'b??11 : new_n850_ = 1'b1;
default : new_n850_ = 1'b0;
endcase
casez ({new_n2746_, new_n1145_})
2'b1? : new_n851_ = 1'b1;
2'b?1 : new_n851_ = 1'b1;
default : new_n851_ = 1'b0;
endcase
casez ({new_n118_, new_n221_, new_n162_, new_n247_})
4'b11?? : new_n852_ = 1'b1;
4'b??11 : new_n852_ = 1'b1;
default : new_n852_ = 1'b0;
endcase
casez ({new_n1632_, new_n1906_})
2'b1? : new_n853_ = 1'b1;
2'b?1 : new_n853_ = 1'b1;
default : new_n853_ = 1'b0;
endcase
casez ({new_n131_, new_n155_})
2'b11 : new_n854_ = 1'b1;
default : new_n854_ = 1'b0;
endcase
casez ({x[0], new_n163_})
2'b11 : new_n855_ = 1'b1;
default : new_n855_ = 1'b0;
endcase
casez ({new_n127_, new_n293_})
2'b11 : new_n856_ = 1'b1;
default : new_n856_ = 1'b0;
endcase
casez ({new_n139_, new_n177_})
2'b11 : new_n857_ = 1'b1;
default : new_n857_ = 1'b0;
endcase
casez ({new_n200_, new_n316_})
2'b11 : new_n858_ = 1'b1;
default : new_n858_ = 1'b0;
endcase
casez ({new_n118_, new_n183_})
2'b11 : new_n859_ = 1'b1;
default : new_n859_ = 1'b0;
endcase
casez ({new_n169_, new_n337_})
2'b11 : new_n860_ = 1'b1;
default : new_n860_ = 1'b0;
endcase
casez ({new_n129_, new_n162_})
2'b11 : new_n861_ = 1'b1;
default : new_n861_ = 1'b0;
endcase
casez ({new_n139_, new_n204_})
2'b11 : new_n862_ = 1'b1;
default : new_n862_ = 1'b0;
endcase
casez ({x[2], new_n212_})
2'b01 : new_n863_ = 1'b1;
default : new_n863_ = 1'b0;
endcase
casez ({new_n96_, new_n221_})
2'b11 : new_n864_ = 1'b1;
default : new_n864_ = 1'b0;
endcase
casez ({new_n127_, new_n229_})
2'b11 : new_n865_ = 1'b1;
default : new_n865_ = 1'b0;
endcase
casez ({new_n142_, new_n231_})
2'b11 : new_n866_ = 1'b1;
default : new_n866_ = 1'b0;
endcase
casez ({new_n124_, new_n136_})
2'b11 : new_n867_ = 1'b1;
default : new_n867_ = 1'b0;
endcase
casez ({new_n97_, new_n143_})
2'b11 : new_n868_ = 1'b1;
default : new_n868_ = 1'b0;
endcase
casez ({x[1], new_n151_})
2'b01 : new_n869_ = 1'b1;
default : new_n869_ = 1'b0;
endcase
casez ({new_n87_, new_n156_})
2'b01 : new_n870_ = 1'b1;
default : new_n870_ = 1'b0;
endcase
casez ({x[1], new_n176_})
2'b01 : new_n871_ = 1'b1;
default : new_n871_ = 1'b0;
endcase
casez ({u[2], new_n191_})
2'b11 : new_n872_ = 1'b1;
default : new_n872_ = 1'b0;
endcase
casez ({u[0], new_n119_})
2'b11 : new_n873_ = 1'b1;
default : new_n873_ = 1'b0;
endcase
casez ({new_n98_, new_n116_})
2'b11 : new_n874_ = 1'b1;
default : new_n874_ = 1'b0;
endcase
casez ({u[0], new_n126_})
2'b11 : new_n875_ = 1'b1;
default : new_n875_ = 1'b0;
endcase
casez ({new_n118_, new_n157_, new_n2128_})
3'b11? : new_n876_ = 1'b1;
3'b??1 : new_n876_ = 1'b1;
default : new_n876_ = 1'b0;
endcase
casez ({new_n311_, new_n618_})
2'b00 : new_n877_ = 1'b1;
default : new_n877_ = 1'b0;
endcase
casez ({new_n93_, new_n272_, new_n175_, new_n211_})
4'b11?? : new_n878_ = 1'b1;
4'b??11 : new_n878_ = 1'b1;
default : new_n878_ = 1'b0;
endcase
casez ({new_n115_, new_n483_, new_n131_, new_n555_})
4'b11?? : new_n879_ = 1'b1;
4'b??11 : new_n879_ = 1'b1;
default : new_n879_ = 1'b0;
endcase
casez ({new_n2116_, new_n131_, new_n144_})
3'b1?? : new_n880_ = 1'b1;
3'b?11 : new_n880_ = 1'b1;
default : new_n880_ = 1'b0;
endcase
casez ({new_n1717_, new_n2117_})
2'b1? : new_n881_ = 1'b1;
2'b?1 : new_n881_ = 1'b1;
default : new_n881_ = 1'b0;
endcase
casez ({new_n96_, new_n295_, new_n3549_})
3'b11? : new_n882_ = 1'b1;
3'b??1 : new_n882_ = 1'b1;
default : new_n882_ = 1'b0;
endcase
casez ({new_n505_, new_n578_})
2'b00 : new_n883_ = 1'b1;
default : new_n883_ = 1'b0;
endcase
casez ({new_n2821_, new_n95_, new_n582_})
3'b1?? : new_n884_ = 1'b1;
3'b?11 : new_n884_ = 1'b1;
default : new_n884_ = 1'b0;
endcase
casez ({new_n2125_, new_n2682_})
2'b1? : new_n885_ = 1'b1;
2'b?1 : new_n885_ = 1'b1;
default : new_n885_ = 1'b0;
endcase
casez ({x[1], new_n244_, new_n599_, new_n580_})
4'b011? : new_n886_ = 1'b1;
4'b???1 : new_n886_ = 1'b1;
default : new_n886_ = 1'b0;
endcase
casez ({new_n138_, new_n553_, new_n160_, new_n600_})
4'b11?? : new_n887_ = 1'b1;
4'b??11 : new_n887_ = 1'b1;
default : new_n887_ = 1'b0;
endcase
casez ({new_n219_, new_n353_, new_n241_, new_n378_})
4'b11?? : new_n888_ = 1'b1;
4'b??11 : new_n888_ = 1'b1;
default : new_n888_ = 1'b0;
endcase
casez ({new_n150_, new_n175_, new_n2830_})
3'b11? : new_n889_ = 1'b1;
3'b??1 : new_n889_ = 1'b1;
default : new_n889_ = 1'b0;
endcase
casez ({new_n1479_, new_n1130_})
2'b1? : new_n890_ = 1'b1;
2'b?1 : new_n890_ = 1'b1;
default : new_n890_ = 1'b0;
endcase
casez ({new_n1347_, new_n1482_})
2'b1? : new_n891_ = 1'b1;
2'b?1 : new_n891_ = 1'b1;
default : new_n891_ = 1'b0;
endcase
casez ({v[2], new_n395_, new_n82_, new_n251_})
4'b01?? : new_n892_ = 1'b1;
4'b??11 : new_n892_ = 1'b1;
default : new_n892_ = 1'b0;
endcase
casez ({new_n89_, new_n404_, new_n118_, new_n199_})
4'b11?? : new_n893_ = 1'b1;
4'b??11 : new_n893_ = 1'b1;
default : new_n893_ = 1'b0;
endcase
casez ({new_n1501_, new_n281_, new_n417_})
3'b1?? : new_n894_ = 1'b1;
3'b?11 : new_n894_ = 1'b1;
default : new_n894_ = 1'b0;
endcase
casez ({new_n2155_, new_n1741_})
2'b1? : new_n895_ = 1'b1;
2'b?1 : new_n895_ = 1'b1;
default : new_n895_ = 1'b0;
endcase
casez ({new_n4664_, new_n139_, new_n191_})
3'b1?? : new_n896_ = 1'b1;
3'b?11 : new_n896_ = 1'b1;
default : new_n896_ = 1'b0;
endcase
casez ({new_n84_, new_n122_})
2'b11 : new_n897_ = 1'b1;
default : new_n897_ = 1'b0;
endcase
casez ({new_n105_, new_n141_})
2'b11 : new_n898_ = 1'b1;
default : new_n898_ = 1'b0;
endcase
casez ({new_n84_, new_n265_})
2'b11 : new_n899_ = 1'b1;
default : new_n899_ = 1'b0;
endcase
casez ({u[0], new_n543_})
2'b01 : new_n900_ = 1'b1;
default : new_n900_ = 1'b0;
endcase
casez ({y[2], new_n292_})
2'b11 : new_n901_ = 1'b1;
default : new_n901_ = 1'b0;
endcase
casez ({new_n110_, new_n169_})
2'b11 : new_n902_ = 1'b1;
default : new_n902_ = 1'b0;
endcase
casez ({new_n154_, new_n186_})
2'b11 : new_n903_ = 1'b1;
default : new_n903_ = 1'b0;
endcase
casez ({new_n104_, new_n339_})
2'b11 : new_n904_ = 1'b1;
default : new_n904_ = 1'b0;
endcase
casez ({x[0], new_n345_})
2'b01 : new_n905_ = 1'b1;
default : new_n905_ = 1'b0;
endcase
casez ({new_n88_, new_n348_})
2'b10 : new_n906_ = 1'b1;
default : new_n906_ = 1'b0;
endcase
casez ({new_n104_, new_n371_})
2'b11 : new_n907_ = 1'b1;
default : new_n907_ = 1'b0;
endcase
casez ({new_n86_, new_n372_})
2'b11 : new_n908_ = 1'b1;
default : new_n908_ = 1'b0;
endcase
casez ({new_n110_, new_n214_})
2'b11 : new_n909_ = 1'b1;
default : new_n909_ = 1'b0;
endcase
casez ({new_n92_, new_n245_})
2'b11 : new_n910_ = 1'b1;
default : new_n910_ = 1'b0;
endcase
casez ({new_n419_, new_n544_})
2'b00 : new_n911_ = 1'b1;
default : new_n911_ = 1'b0;
endcase
casez ({y[2], new_n164_, new_n1525_})
3'b11? : new_n912_ = 1'b1;
3'b??1 : new_n912_ = 1'b1;
default : new_n912_ = 1'b0;
endcase
casez ({v[2], new_n292_, new_n82_, new_n277_})
4'b01?? : new_n913_ = 1'b1;
4'b??01 : new_n913_ = 1'b1;
default : new_n913_ = 1'b0;
endcase
casez ({new_n139_, new_n168_, new_n150_, new_n164_})
4'b11?? : new_n914_ = 1'b1;
4'b??11 : new_n914_ = 1'b1;
default : new_n914_ = 1'b0;
endcase
casez ({new_n79_, new_n269_})
2'b11 : new_n915_ = 1'b1;
default : new_n915_ = 1'b0;
endcase
casez ({y[2], new_n277_})
2'b11 : new_n916_ = 1'b1;
default : new_n916_ = 1'b0;
endcase
casez ({y[2], new_n283_})
2'b11 : new_n917_ = 1'b1;
default : new_n917_ = 1'b0;
endcase
casez ({new_n353_, new_n1942_, new_n736_})
3'b11? : new_n918_ = 1'b1;
3'b??1 : new_n918_ = 1'b1;
default : new_n918_ = 1'b0;
endcase
casez ({new_n373_, new_n739_, new_n438_, new_n562_})
4'b11?? : new_n919_ = 1'b1;
4'b??11 : new_n919_ = 1'b1;
default : new_n919_ = 1'b0;
endcase
casez ({new_n4616_, new_n913_})
2'b1? : new_n920_ = 1'b1;
2'b?1 : new_n920_ = 1'b1;
default : new_n920_ = 1'b0;
endcase
casez ({new_n82_, new_n698_, new_n104_, new_n626_})
4'b11?? : new_n921_ = 1'b1;
4'b??11 : new_n921_ = 1'b1;
default : new_n921_ = 1'b0;
endcase
casez ({new_n331_, new_n1808_, new_n921_})
3'b11? : new_n922_ = 1'b1;
3'b??1 : new_n922_ = 1'b1;
default : new_n922_ = 1'b0;
endcase
casez ({x[1], v[1]})
2'b10 : new_n923_ = 1'b1;
default : new_n923_ = 1'b0;
endcase
casez ({y[1], v[0]})
2'b01 : new_n924_ = 1'b1;
default : new_n924_ = 1'b0;
endcase
casez ({new_n89_, new_n101_})
2'b00 : new_n925_ = 1'b1;
default : new_n925_ = 1'b0;
endcase
casez ({x[0], new_n86_})
2'b10 : new_n926_ = 1'b1;
default : new_n926_ = 1'b0;
endcase
casez ({y[1], new_n91_})
2'b11 : new_n927_ = 1'b1;
default : new_n927_ = 1'b0;
endcase
casez ({new_n166_, new_n174_})
2'b00 : new_n928_ = 1'b1;
default : new_n928_ = 1'b0;
endcase
casez ({new_n3398_, new_n3389_})
2'b1? : new_n929_ = 1'b1;
2'b?1 : new_n929_ = 1'b1;
default : new_n929_ = 1'b0;
endcase
casez ({new_n158_, new_n251_})
2'b00 : new_n930_ = 1'b1;
default : new_n930_ = 1'b0;
endcase
casez ({new_n251_, new_n254_})
2'b00 : new_n931_ = 1'b1;
default : new_n931_ = 1'b0;
endcase
casez ({new_n1110_, new_n237_})
2'b1? : new_n932_ = 1'b1;
2'b?1 : new_n932_ = 1'b1;
default : new_n932_ = 1'b0;
endcase
casez ({new_n161_, new_n166_})
2'b00 : new_n933_ = 1'b1;
default : new_n933_ = 1'b0;
endcase
casez ({new_n159_, new_n170_})
2'b00 : new_n934_ = 1'b1;
default : new_n934_ = 1'b0;
endcase
casez ({new_n183_, new_n347_})
2'b00 : new_n935_ = 1'b1;
default : new_n935_ = 1'b0;
endcase
casez ({new_n196_, new_n204_})
2'b00 : new_n936_ = 1'b1;
default : new_n936_ = 1'b0;
endcase
casez ({new_n124_, new_n141_})
2'b11 : new_n937_ = 1'b1;
default : new_n937_ = 1'b0;
endcase
casez ({new_n127_, new_n153_})
2'b11 : new_n938_ = 1'b1;
default : new_n938_ = 1'b0;
endcase
casez ({new_n131_, new_n300_})
2'b11 : new_n939_ = 1'b1;
default : new_n939_ = 1'b0;
endcase
casez ({x[0], new_n163_})
2'b01 : new_n940_ = 1'b1;
default : new_n940_ = 1'b0;
endcase
casez ({new_n139_, new_n158_})
2'b11 : new_n941_ = 1'b1;
default : new_n941_ = 1'b0;
endcase
casez ({new_n127_, new_n169_})
2'b11 : new_n942_ = 1'b1;
default : new_n942_ = 1'b0;
endcase
casez ({new_n80_, new_n177_})
2'b01 : new_n943_ = 1'b1;
default : new_n943_ = 1'b0;
endcase
casez ({new_n150_, new_n177_})
2'b11 : new_n944_ = 1'b1;
default : new_n944_ = 1'b0;
endcase
casez ({new_n226_, new_n332_})
2'b11 : new_n945_ = 1'b1;
default : new_n945_ = 1'b0;
endcase
casez ({new_n150_, new_n192_})
2'b11 : new_n946_ = 1'b1;
default : new_n946_ = 1'b0;
endcase
casez ({new_n150_, new_n210_})
2'b11 : new_n947_ = 1'b1;
default : new_n947_ = 1'b0;
endcase
casez ({new_n158_, new_n211_})
2'b11 : new_n948_ = 1'b1;
default : new_n948_ = 1'b0;
endcase
casez ({new_n127_, new_n237_})
2'b11 : new_n949_ = 1'b1;
default : new_n949_ = 1'b0;
endcase
casez ({new_n107_, new_n133_})
2'b01 : new_n950_ = 1'b1;
default : new_n950_ = 1'b0;
endcase
casez ({new_n220_, new_n248_})
2'b11 : new_n951_ = 1'b1;
default : new_n951_ = 1'b0;
endcase
casez ({y[2], new_n126_})
2'b01 : new_n952_ = 1'b1;
default : new_n952_ = 1'b0;
endcase
casez ({new_n82_, new_n147_})
2'b01 : new_n953_ = 1'b1;
default : new_n953_ = 1'b0;
endcase
casez ({new_n138_, new_n148_})
2'b11 : new_n954_ = 1'b1;
default : new_n954_ = 1'b0;
endcase
casez ({y[2], new_n173_})
2'b01 : new_n955_ = 1'b1;
default : new_n955_ = 1'b0;
endcase
casez ({u[2], new_n196_})
2'b11 : new_n956_ = 1'b1;
default : new_n956_ = 1'b0;
endcase
casez ({x[2], new_n148_})
2'b11 : new_n957_ = 1'b1;
default : new_n957_ = 1'b0;
endcase
casez ({new_n98_, new_n126_})
2'b11 : new_n958_ = 1'b1;
default : new_n958_ = 1'b0;
endcase
casez ({v[1], new_n123_})
2'b11 : new_n959_ = 1'b1;
default : new_n959_ = 1'b0;
endcase
casez ({v[1], new_n123_})
2'b01 : new_n960_ = 1'b1;
default : new_n960_ = 1'b0;
endcase
casez ({new_n79_, new_n128_})
2'b11 : new_n961_ = 1'b1;
default : new_n961_ = 1'b0;
endcase
casez ({v[1], new_n129_})
2'b01 : new_n962_ = 1'b1;
default : new_n962_ = 1'b0;
endcase
casez ({u[1], new_n131_})
2'b01 : new_n963_ = 1'b1;
default : new_n963_ = 1'b0;
endcase
casez ({x[0], new_n135_})
2'b11 : new_n964_ = 1'b1;
default : new_n964_ = 1'b0;
endcase
casez ({new_n86_, new_n115_})
2'b11 : new_n965_ = 1'b1;
default : new_n965_ = 1'b0;
endcase
casez ({new_n360_, new_n480_})
2'b00 : new_n966_ = 1'b1;
default : new_n966_ = 1'b0;
endcase
casez ({new_n3588_, new_n286_})
2'b1? : new_n967_ = 1'b1;
2'b?1 : new_n967_ = 1'b1;
default : new_n967_ = 1'b0;
endcase
casez ({new_n323_, new_n607_})
2'b00 : new_n968_ = 1'b1;
default : new_n968_ = 1'b0;
endcase
casez ({new_n106_, new_n360_})
2'b00 : new_n969_ = 1'b1;
default : new_n969_ = 1'b0;
endcase
casez ({new_n1642_, new_n682_})
2'b1? : new_n970_ = 1'b1;
2'b?1 : new_n970_ = 1'b1;
default : new_n970_ = 1'b0;
endcase
casez ({new_n295_, new_n423_})
2'b00 : new_n971_ = 1'b1;
default : new_n971_ = 1'b0;
endcase
casez ({new_n245_, new_n450_})
2'b00 : new_n972_ = 1'b1;
default : new_n972_ = 1'b0;
endcase
casez ({u[0], new_n295_})
2'b01 : new_n973_ = 1'b1;
default : new_n973_ = 1'b0;
endcase
casez ({x[0], new_n579_})
2'b01 : new_n974_ = 1'b1;
default : new_n974_ = 1'b0;
endcase
casez ({new_n94_, new_n329_})
2'b11 : new_n975_ = 1'b1;
default : new_n975_ = 1'b0;
endcase
casez ({y[0], new_n681_})
2'b11 : new_n976_ = 1'b1;
default : new_n976_ = 1'b0;
endcase
casez ({new_n114_, new_n133_})
2'b11 : new_n977_ = 1'b1;
default : new_n977_ = 1'b0;
endcase
casez ({new_n110_, new_n250_})
2'b11 : new_n978_ = 1'b1;
default : new_n978_ = 1'b0;
endcase
casez ({new_n83_, new_n267_})
2'b11 : new_n979_ = 1'b1;
default : new_n979_ = 1'b0;
endcase
casez ({new_n103_, new_n271_})
2'b11 : new_n980_ = 1'b1;
default : new_n980_ = 1'b0;
endcase
casez ({new_n131_, new_n157_})
2'b11 : new_n981_ = 1'b1;
default : new_n981_ = 1'b0;
endcase
casez ({x[0], new_n157_})
2'b01 : new_n982_ = 1'b1;
default : new_n982_ = 1'b0;
endcase
casez ({u[0], new_n282_})
2'b01 : new_n983_ = 1'b1;
default : new_n983_ = 1'b0;
endcase
casez ({v[1], new_n175_})
2'b11 : new_n984_ = 1'b1;
default : new_n984_ = 1'b0;
endcase
casez ({new_n80_, new_n325_})
2'b11 : new_n985_ = 1'b1;
default : new_n985_ = 1'b0;
endcase
casez ({new_n103_, new_n330_})
2'b11 : new_n986_ = 1'b1;
default : new_n986_ = 1'b0;
endcase
casez ({u[0], new_n225_})
2'b11 : new_n987_ = 1'b1;
default : new_n987_ = 1'b0;
endcase
casez ({new_n121_, new_n139_})
2'b11 : new_n988_ = 1'b1;
default : new_n988_ = 1'b0;
endcase
casez ({new_n195_, new_n674_})
2'b00 : new_n989_ = 1'b1;
default : new_n989_ = 1'b0;
endcase
casez ({u[0], new_n168_})
2'b11 : new_n990_ = 1'b1;
default : new_n990_ = 1'b0;
endcase
casez ({x[0], x[1]})
2'b00 : new_n991_ = 1'b1;
default : new_n991_ = 1'b0;
endcase
casez ({new_n85_, new_n305_})
2'b00 : new_n992_ = 1'b1;
default : new_n992_ = 1'b0;
endcase
casez ({new_n224_, new_n284_})
2'b00 : new_n993_ = 1'b1;
default : new_n993_ = 1'b0;
endcase
casez ({new_n234_, new_n257_})
2'b11 : new_n994_ = 1'b1;
default : new_n994_ = 1'b0;
endcase
casez ({new_n3455_, new_n251_})
2'b1? : new_n995_ = 1'b1;
2'b?1 : new_n995_ = 1'b1;
default : new_n995_ = 1'b0;
endcase
casez ({u[2], new_n242_, new_n293_})
3'b01? : new_n996_ = 1'b1;
3'b??1 : new_n996_ = 1'b1;
default : new_n996_ = 1'b0;
endcase
casez ({new_n1363_, new_n183_})
2'b1? : new_n997_ = 1'b1;
2'b?1 : new_n997_ = 1'b1;
default : new_n997_ = 1'b0;
endcase
casez ({new_n129_, new_n221_})
2'b00 : new_n998_ = 1'b1;
default : new_n998_ = 1'b0;
endcase
casez ({new_n94_, new_n228_})
2'b00 : new_n999_ = 1'b1;
default : new_n999_ = 1'b0;
endcase
casez ({new_n208_, new_n242_})
2'b00 : new_n1000_ = 1'b1;
default : new_n1000_ = 1'b0;
endcase
casez ({new_n82_, new_n141_})
2'b01 : new_n1001_ = 1'b1;
default : new_n1001_ = 1'b0;
endcase
casez ({new_n83_, new_n140_})
2'b01 : new_n1002_ = 1'b1;
default : new_n1002_ = 1'b0;
endcase
casez ({new_n229_, new_n260_})
2'b11 : new_n1003_ = 1'b1;
default : new_n1003_ = 1'b0;
endcase
casez ({new_n169_, new_n261_})
2'b11 : new_n1004_ = 1'b1;
default : new_n1004_ = 1'b0;
endcase
casez ({new_n124_, new_n146_})
2'b11 : new_n1005_ = 1'b1;
default : new_n1005_ = 1'b0;
endcase
casez ({y[2], new_n1005_, new_n216_, new_n542_})
4'b11?? : new_n1006_ = 1'b1;
4'b??11 : new_n1006_ = 1'b1;
default : new_n1006_ = 1'b0;
endcase
casez ({new_n123_, new_n148_})
2'b11 : new_n1007_ = 1'b1;
default : new_n1007_ = 1'b0;
endcase
casez ({new_n138_, new_n273_})
2'b11 : new_n1008_ = 1'b1;
default : new_n1008_ = 1'b0;
endcase
casez ({new_n118_, new_n159_})
2'b11 : new_n1009_ = 1'b1;
default : new_n1009_ = 1'b0;
endcase
casez ({new_n150_, new_n160_})
2'b11 : new_n1010_ = 1'b1;
default : new_n1010_ = 1'b0;
endcase
casez ({new_n140_, new_n162_})
2'b11 : new_n1011_ = 1'b1;
default : new_n1011_ = 1'b0;
endcase
casez ({new_n115_, new_n161_})
2'b11 : new_n1012_ = 1'b1;
default : new_n1012_ = 1'b0;
endcase
casez ({v[2], new_n165_})
2'b01 : new_n1013_ = 1'b1;
default : new_n1013_ = 1'b0;
endcase
casez ({new_n131_, new_n166_})
2'b11 : new_n1014_ = 1'b1;
default : new_n1014_ = 1'b0;
endcase
casez ({new_n150_, new_n167_})
2'b11 : new_n1015_ = 1'b1;
default : new_n1015_ = 1'b0;
endcase
casez ({new_n79_, new_n170_})
2'b01 : new_n1016_ = 1'b1;
default : new_n1016_ = 1'b0;
endcase
casez ({new_n201_, new_n316_})
2'b11 : new_n1017_ = 1'b1;
default : new_n1017_ = 1'b0;
endcase
casez ({new_n162_, new_n173_})
2'b11 : new_n1018_ = 1'b1;
default : new_n1018_ = 1'b0;
endcase
casez ({v[1], new_n189_})
2'b11 : new_n1019_ = 1'b1;
default : new_n1019_ = 1'b0;
endcase
casez ({x[1], new_n196_})
2'b01 : new_n1020_ = 1'b1;
default : new_n1020_ = 1'b0;
endcase
casez ({new_n115_, new_n151_})
2'b11 : new_n1021_ = 1'b1;
default : new_n1021_ = 1'b0;
endcase
casez ({new_n161_, new_n358_})
2'b11 : new_n1022_ = 1'b1;
default : new_n1022_ = 1'b0;
endcase
casez ({new_n80_, new_n204_})
2'b01 : new_n1023_ = 1'b1;
default : new_n1023_ = 1'b0;
endcase
casez ({new_n80_, new_n206_})
2'b01 : new_n1024_ = 1'b1;
default : new_n1024_ = 1'b0;
endcase
casez ({new_n101_, new_n207_})
2'b11 : new_n1025_ = 1'b1;
default : new_n1025_ = 1'b0;
endcase
casez ({new_n160_, new_n369_})
2'b11 : new_n1026_ = 1'b1;
default : new_n1026_ = 1'b0;
endcase
casez ({new_n177_, new_n211_})
2'b11 : new_n1027_ = 1'b1;
default : new_n1027_ = 1'b0;
endcase
casez ({new_n104_, new_n211_})
2'b11 : new_n1028_ = 1'b1;
default : new_n1028_ = 1'b0;
endcase
casez ({x[1], new_n206_})
2'b11 : new_n1029_ = 1'b1;
default : new_n1029_ = 1'b0;
endcase
casez ({new_n127_, new_n212_})
2'b11 : new_n1030_ = 1'b1;
default : new_n1030_ = 1'b0;
endcase
casez ({new_n97_, new_n222_})
2'b11 : new_n1031_ = 1'b1;
default : new_n1031_ = 1'b0;
endcase
casez ({new_n194_, new_n244_})
2'b11 : new_n1032_ = 1'b1;
default : new_n1032_ = 1'b0;
endcase
casez ({new_n261_, new_n660_, new_n766_, new_n1032_})
4'b11?? : new_n1033_ = 1'b1;
4'b??11 : new_n1033_ = 1'b1;
default : new_n1033_ = 1'b0;
endcase
casez ({v[2], new_n136_})
2'b11 : new_n1034_ = 1'b1;
default : new_n1034_ = 1'b0;
endcase
casez ({y[1], new_n136_})
2'b01 : new_n1035_ = 1'b1;
default : new_n1035_ = 1'b0;
endcase
casez ({new_n95_, new_n248_})
2'b11 : new_n1036_ = 1'b1;
default : new_n1036_ = 1'b0;
endcase
casez ({new_n137_, new_n250_})
2'b11 : new_n1037_ = 1'b1;
default : new_n1037_ = 1'b0;
endcase
casez ({new_n84_, new_n145_})
2'b11 : new_n1038_ = 1'b1;
default : new_n1038_ = 1'b0;
endcase
casez ({new_n79_, new_n151_})
2'b01 : new_n1039_ = 1'b1;
default : new_n1039_ = 1'b0;
endcase
casez ({x[1], new_n167_})
2'b11 : new_n1040_ = 1'b1;
default : new_n1040_ = 1'b0;
endcase
casez ({v[1], new_n189_})
2'b01 : new_n1041_ = 1'b1;
default : new_n1041_ = 1'b0;
endcase
casez ({u[2], new_n201_})
2'b11 : new_n1042_ = 1'b1;
default : new_n1042_ = 1'b0;
endcase
casez ({new_n131_, new_n401_})
2'b11 : new_n1043_ = 1'b1;
default : new_n1043_ = 1'b0;
endcase
casez ({new_n95_, new_n115_})
2'b11 : new_n1044_ = 1'b1;
default : new_n1044_ = 1'b0;
endcase
casez ({new_n89_, new_n124_})
2'b11 : new_n1045_ = 1'b1;
default : new_n1045_ = 1'b0;
endcase
casez ({new_n104_, new_n139_})
2'b11 : new_n1046_ = 1'b1;
default : new_n1046_ = 1'b0;
endcase
casez ({x[2], new_n131_})
2'b11 : new_n1047_ = 1'b1;
default : new_n1047_ = 1'b0;
endcase
casez ({new_n2145_, new_n779_})
2'b1? : new_n1048_ = 1'b1;
2'b?1 : new_n1048_ = 1'b1;
default : new_n1048_ = 1'b0;
endcase
casez ({new_n1798_, new_n271_})
2'b1? : new_n1049_ = 1'b1;
2'b?1 : new_n1049_ = 1'b1;
default : new_n1049_ = 1'b0;
endcase
casez ({new_n1609_, new_n367_})
2'b1? : new_n1050_ = 1'b1;
2'b?1 : new_n1050_ = 1'b1;
default : new_n1050_ = 1'b0;
endcase
casez ({new_n137_, new_n214_, new_n668_})
3'b11? : new_n1051_ = 1'b1;
3'b??1 : new_n1051_ = 1'b1;
default : new_n1051_ = 1'b0;
endcase
casez ({new_n83_, new_n226_, new_n683_})
3'b11? : new_n1052_ = 1'b1;
3'b??1 : new_n1052_ = 1'b1;
default : new_n1052_ = 1'b0;
endcase
casez ({new_n245_, new_n442_})
2'b00 : new_n1053_ = 1'b1;
default : new_n1053_ = 1'b0;
endcase
casez ({new_n92_, new_n253_})
2'b11 : new_n1054_ = 1'b1;
default : new_n1054_ = 1'b0;
endcase
casez ({new_n80_, new_n259_})
2'b11 : new_n1055_ = 1'b1;
default : new_n1055_ = 1'b0;
endcase
casez ({new_n157_, new_n273_})
2'b11 : new_n1056_ = 1'b1;
default : new_n1056_ = 1'b0;
endcase
casez ({v[1], new_n292_})
2'b01 : new_n1057_ = 1'b1;
default : new_n1057_ = 1'b0;
endcase
casez ({u[0], new_n294_})
2'b01 : new_n1058_ = 1'b1;
default : new_n1058_ = 1'b0;
endcase
casez ({x[0], new_n294_})
2'b11 : new_n1059_ = 1'b1;
default : new_n1059_ = 1'b0;
endcase
casez ({new_n112_, new_n169_})
2'b11 : new_n1060_ = 1'b1;
default : new_n1060_ = 1'b0;
endcase
casez ({new_n94_, new_n308_})
2'b11 : new_n1061_ = 1'b1;
default : new_n1061_ = 1'b0;
endcase
casez ({v[2], new_n308_})
2'b01 : new_n1062_ = 1'b1;
default : new_n1062_ = 1'b0;
endcase
casez ({new_n81_, new_n329_})
2'b11 : new_n1063_ = 1'b1;
default : new_n1063_ = 1'b0;
endcase
casez ({new_n104_, new_n330_})
2'b11 : new_n1064_ = 1'b1;
default : new_n1064_ = 1'b0;
endcase
casez ({new_n104_, new_n378_})
2'b11 : new_n1065_ = 1'b1;
default : new_n1065_ = 1'b0;
endcase
casez ({new_n85_, new_n387_})
2'b11 : new_n1066_ = 1'b1;
default : new_n1066_ = 1'b0;
endcase
casez ({new_n81_, new_n395_})
2'b11 : new_n1067_ = 1'b1;
default : new_n1067_ = 1'b0;
endcase
casez ({y[0], new_n408_})
2'b01 : new_n1068_ = 1'b1;
default : new_n1068_ = 1'b0;
endcase
casez ({new_n88_, new_n455_})
2'b11 : new_n1069_ = 1'b1;
default : new_n1069_ = 1'b0;
endcase
casez ({new_n115_, new_n175_})
2'b11 : new_n1070_ = 1'b1;
default : new_n1070_ = 1'b0;
endcase
casez ({v[1], new_n186_})
2'b01 : new_n1071_ = 1'b1;
default : new_n1071_ = 1'b0;
endcase
casez ({new_n157_, new_n198_})
2'b11 : new_n1072_ = 1'b1;
default : new_n1072_ = 1'b0;
endcase
casez ({new_n89_, new_n122_})
2'b11 : new_n1073_ = 1'b1;
default : new_n1073_ = 1'b0;
endcase
casez ({new_n1945_, new_n188_})
2'b1? : new_n1074_ = 1'b1;
2'b?1 : new_n1074_ = 1'b1;
default : new_n1074_ = 1'b0;
endcase
casez ({new_n2742_, new_n368_})
2'b1? : new_n1075_ = 1'b1;
2'b?1 : new_n1075_ = 1'b1;
default : new_n1075_ = 1'b0;
endcase
casez ({new_n2835_, new_n312_})
2'b1? : new_n1076_ = 1'b1;
2'b?1 : new_n1076_ = 1'b1;
default : new_n1076_ = 1'b0;
endcase
casez ({new_n2750_, new_n575_})
2'b1? : new_n1077_ = 1'b1;
2'b?1 : new_n1077_ = 1'b1;
default : new_n1077_ = 1'b0;
endcase
casez ({new_n162_, new_n235_, new_n610_})
3'b11? : new_n1078_ = 1'b1;
3'b??1 : new_n1078_ = 1'b1;
default : new_n1078_ = 1'b0;
endcase
casez ({new_n2832_, new_n613_})
2'b1? : new_n1079_ = 1'b1;
2'b?1 : new_n1079_ = 1'b1;
default : new_n1079_ = 1'b0;
endcase
casez ({new_n2849_, new_n617_})
2'b1? : new_n1080_ = 1'b1;
2'b?1 : new_n1080_ = 1'b1;
default : new_n1080_ = 1'b0;
endcase
casez ({new_n127_, new_n317_, new_n625_})
3'b11? : new_n1081_ = 1'b1;
3'b??1 : new_n1081_ = 1'b1;
default : new_n1081_ = 1'b0;
endcase
casez ({new_n312_, new_n637_})
2'b00 : new_n1082_ = 1'b1;
default : new_n1082_ = 1'b0;
endcase
casez ({new_n173_, new_n273_, new_n655_})
3'b11? : new_n1083_ = 1'b1;
3'b??1 : new_n1083_ = 1'b1;
default : new_n1083_ = 1'b0;
endcase
casez ({new_n281_, new_n338_, new_n402_})
3'b11? : new_n1084_ = 1'b1;
3'b??1 : new_n1084_ = 1'b1;
default : new_n1084_ = 1'b0;
endcase
casez ({y[1], new_n750_, new_n464_})
3'b11? : new_n1085_ = 1'b1;
3'b??1 : new_n1085_ = 1'b1;
default : new_n1085_ = 1'b0;
endcase
casez ({new_n3463_, new_n477_})
2'b1? : new_n1086_ = 1'b1;
2'b?1 : new_n1086_ = 1'b1;
default : new_n1086_ = 1'b0;
endcase
casez ({new_n84_, new_n263_})
2'b11 : new_n1087_ = 1'b1;
default : new_n1087_ = 1'b0;
endcase
casez ({new_n117_, new_n214_})
2'b11 : new_n1088_ = 1'b1;
default : new_n1088_ = 1'b0;
endcase
casez ({y[2], new_n331_})
2'b01 : new_n1089_ = 1'b1;
default : new_n1089_ = 1'b0;
endcase
casez ({v[0], v[1]})
2'b00 : new_n1090_ = 1'b1;
default : new_n1090_ = 1'b0;
endcase
casez ({new_n88_, new_n346_})
2'b00 : new_n1091_ = 1'b1;
default : new_n1091_ = 1'b0;
endcase
casez ({u[2], new_n103_})
2'b01 : new_n1092_ = 1'b1;
default : new_n1092_ = 1'b0;
endcase
casez ({y[0], new_n82_})
2'b00 : new_n1093_ = 1'b1;
default : new_n1093_ = 1'b0;
endcase
casez ({new_n80_, new_n85_})
2'b01 : new_n1094_ = 1'b1;
default : new_n1094_ = 1'b0;
endcase
casez ({new_n86_, new_n88_})
2'b01 : new_n1095_ = 1'b1;
default : new_n1095_ = 1'b0;
endcase
casez ({new_n82_, new_n90_})
2'b01 : new_n1096_ = 1'b1;
default : new_n1096_ = 1'b0;
endcase
casez ({new_n86_, new_n96_})
2'b01 : new_n1097_ = 1'b1;
default : new_n1097_ = 1'b0;
endcase
casez ({new_n80_, new_n242_})
2'b01 : new_n1098_ = 1'b1;
default : new_n1098_ = 1'b0;
endcase
casez ({new_n89_, new_n94_})
2'b11 : new_n1099_ = 1'b1;
default : new_n1099_ = 1'b0;
endcase
casez ({new_n140_, new_n173_})
2'b00 : new_n1100_ = 1'b1;
default : new_n1100_ = 1'b0;
endcase
casez ({new_n158_, new_n242_})
2'b00 : new_n1101_ = 1'b1;
default : new_n1101_ = 1'b0;
endcase
casez ({new_n84_, new_n140_})
2'b01 : new_n1102_ = 1'b1;
default : new_n1102_ = 1'b0;
endcase
casez ({new_n77_, new_n141_})
2'b11 : new_n1103_ = 1'b1;
default : new_n1103_ = 1'b0;
endcase
casez ({new_n127_, new_n142_})
2'b11 : new_n1104_ = 1'b1;
default : new_n1104_ = 1'b0;
endcase
casez ({new_n235_, new_n257_})
2'b11 : new_n1105_ = 1'b1;
default : new_n1105_ = 1'b0;
endcase
casez ({new_n162_, new_n261_})
2'b11 : new_n1106_ = 1'b1;
default : new_n1106_ = 1'b0;
endcase
casez ({u[1], new_n264_})
2'b01 : new_n1107_ = 1'b1;
default : new_n1107_ = 1'b0;
endcase
casez ({new_n148_, new_n151_})
2'b11 : new_n1108_ = 1'b1;
default : new_n1108_ = 1'b0;
endcase
casez ({new_n129_, new_n153_})
2'b11 : new_n1109_ = 1'b1;
default : new_n1109_ = 1'b0;
endcase
casez ({new_n79_, new_n258_})
2'b01 : new_n1110_ = 1'b1;
default : new_n1110_ = 1'b0;
endcase
casez ({new_n144_, new_n273_})
2'b11 : new_n1111_ = 1'b1;
default : new_n1111_ = 1'b0;
endcase
casez ({new_n118_, new_n158_})
2'b11 : new_n1112_ = 1'b1;
default : new_n1112_ = 1'b0;
endcase
casez ({new_n79_, new_n158_})
2'b11 : new_n1113_ = 1'b1;
default : new_n1113_ = 1'b0;
endcase
casez ({new_n131_, new_n278_})
2'b11 : new_n1114_ = 1'b1;
default : new_n1114_ = 1'b0;
endcase
casez ({new_n139_, new_n278_})
2'b11 : new_n1115_ = 1'b1;
default : new_n1115_ = 1'b0;
endcase
casez ({new_n150_, new_n159_})
2'b11 : new_n1116_ = 1'b1;
default : new_n1116_ = 1'b0;
endcase
casez ({new_n139_, new_n159_})
2'b11 : new_n1117_ = 1'b1;
default : new_n1117_ = 1'b0;
endcase
casez ({new_n115_, new_n160_})
2'b11 : new_n1118_ = 1'b1;
default : new_n1118_ = 1'b0;
endcase
casez ({new_n148_, new_n161_})
2'b11 : new_n1119_ = 1'b1;
default : new_n1119_ = 1'b0;
endcase
casez ({new_n145_, new_n162_})
2'b11 : new_n1120_ = 1'b1;
default : new_n1120_ = 1'b0;
endcase
casez ({new_n118_, new_n166_})
2'b11 : new_n1121_ = 1'b1;
default : new_n1121_ = 1'b0;
endcase
casez ({new_n123_, new_n169_})
2'b11 : new_n1122_ = 1'b1;
default : new_n1122_ = 1'b0;
endcase
casez ({new_n115_, new_n170_})
2'b11 : new_n1123_ = 1'b1;
default : new_n1123_ = 1'b0;
endcase
casez ({new_n118_, new_n300_})
2'b11 : new_n1124_ = 1'b1;
default : new_n1124_ = 1'b0;
endcase
casez ({new_n79_, new_n301_})
2'b01 : new_n1125_ = 1'b1;
default : new_n1125_ = 1'b0;
endcase
casez ({new_n87_, new_n174_})
2'b11 : new_n1126_ = 1'b1;
default : new_n1126_ = 1'b0;
endcase
casez ({new_n194_, new_n306_})
2'b11 : new_n1127_ = 1'b1;
default : new_n1127_ = 1'b0;
endcase
casez ({new_n176_, new_n1127_, new_n372_, new_n790_})
4'b11?? : new_n1128_ = 1'b1;
4'b??11 : new_n1128_ = 1'b1;
default : new_n1128_ = 1'b0;
endcase
casez ({x[1], new_n177_})
2'b11 : new_n1129_ = 1'b1;
default : new_n1129_ = 1'b0;
endcase
casez ({new_n115_, new_n176_})
2'b11 : new_n1130_ = 1'b1;
default : new_n1130_ = 1'b0;
endcase
casez ({new_n131_, new_n183_})
2'b11 : new_n1131_ = 1'b1;
default : new_n1131_ = 1'b0;
endcase
casez ({new_n87_, new_n187_})
2'b01 : new_n1132_ = 1'b1;
default : new_n1132_ = 1'b0;
endcase
casez ({new_n79_, new_n187_})
2'b01 : new_n1133_ = 1'b1;
default : new_n1133_ = 1'b0;
endcase
casez ({x[1], new_n187_})
2'b01 : new_n1134_ = 1'b1;
default : new_n1134_ = 1'b0;
endcase
casez ({y[2], new_n190_})
2'b01 : new_n1135_ = 1'b1;
default : new_n1135_ = 1'b0;
endcase
casez ({new_n150_, new_n196_})
2'b11 : new_n1136_ = 1'b1;
default : new_n1136_ = 1'b0;
endcase
casez ({new_n93_, new_n196_})
2'b01 : new_n1137_ = 1'b1;
default : new_n1137_ = 1'b0;
endcase
casez ({new_n131_, new_n178_})
2'b11 : new_n1138_ = 1'b1;
default : new_n1138_ = 1'b0;
endcase
casez ({new_n161_, new_n209_})
2'b11 : new_n1139_ = 1'b1;
default : new_n1139_ = 1'b0;
endcase
casez ({new_n129_, new_n207_})
2'b11 : new_n1140_ = 1'b1;
default : new_n1140_ = 1'b0;
endcase
casez ({new_n88_, new_n211_})
2'b11 : new_n1141_ = 1'b1;
default : new_n1141_ = 1'b0;
endcase
casez ({new_n103_, new_n211_})
2'b11 : new_n1142_ = 1'b1;
default : new_n1142_ = 1'b0;
endcase
casez ({new_n154_, new_n213_})
2'b11 : new_n1143_ = 1'b1;
default : new_n1143_ = 1'b0;
endcase
casez ({new_n178_, new_n214_})
2'b11 : new_n1144_ = 1'b1;
default : new_n1144_ = 1'b0;
endcase
casez ({new_n200_, new_n216_})
2'b11 : new_n1145_ = 1'b1;
default : new_n1145_ = 1'b0;
endcase
casez ({new_n213_, new_n216_})
2'b11 : new_n1146_ = 1'b1;
default : new_n1146_ = 1'b0;
endcase
casez ({new_n158_, new_n216_})
2'b11 : new_n1147_ = 1'b1;
default : new_n1147_ = 1'b0;
endcase
casez ({new_n154_, new_n221_})
2'b11 : new_n1148_ = 1'b1;
default : new_n1148_ = 1'b0;
endcase
casez ({new_n176_, new_n221_})
2'b11 : new_n1149_ = 1'b1;
default : new_n1149_ = 1'b0;
endcase
casez ({new_n167_, new_n221_})
2'b11 : new_n1150_ = 1'b1;
default : new_n1150_ = 1'b0;
endcase
casez ({new_n118_, new_n224_})
2'b11 : new_n1151_ = 1'b1;
default : new_n1151_ = 1'b0;
endcase
casez ({new_n264_, new_n357_})
2'b11 : new_n1152_ = 1'b1;
default : new_n1152_ = 1'b0;
endcase
casez ({new_n95_, new_n237_})
2'b11 : new_n1153_ = 1'b1;
default : new_n1153_ = 1'b0;
endcase
casez ({new_n229_, new_n244_})
2'b11 : new_n1154_ = 1'b1;
default : new_n1154_ = 1'b0;
endcase
casez ({new_n167_, new_n243_})
2'b11 : new_n1155_ = 1'b1;
default : new_n1155_ = 1'b0;
endcase
casez ({new_n85_, new_n249_})
2'b11 : new_n1156_ = 1'b1;
default : new_n1156_ = 1'b0;
endcase
casez ({new_n127_, new_n251_})
2'b11 : new_n1157_ = 1'b1;
default : new_n1157_ = 1'b0;
endcase
casez ({y[2], new_n140_})
2'b11 : new_n1158_ = 1'b1;
default : new_n1158_ = 1'b0;
endcase
casez ({v[2], new_n141_})
2'b01 : new_n1159_ = 1'b1;
default : new_n1159_ = 1'b0;
endcase
casez ({x[2], new_n142_})
2'b11 : new_n1160_ = 1'b1;
default : new_n1160_ = 1'b0;
endcase
casez ({y[2], new_n144_})
2'b01 : new_n1161_ = 1'b1;
default : new_n1161_ = 1'b0;
endcase
casez ({u[2], new_n158_})
2'b01 : new_n1162_ = 1'b1;
default : new_n1162_ = 1'b0;
endcase
casez ({x[1], new_n159_})
2'b01 : new_n1163_ = 1'b1;
default : new_n1163_ = 1'b0;
endcase
casez ({new_n118_, new_n161_})
2'b11 : new_n1164_ = 1'b1;
default : new_n1164_ = 1'b0;
endcase
casez ({new_n83_, new_n173_})
2'b11 : new_n1165_ = 1'b1;
default : new_n1165_ = 1'b0;
endcase
casez ({new_n81_, new_n180_})
2'b01 : new_n1166_ = 1'b1;
default : new_n1166_ = 1'b0;
endcase
casez ({u[2], new_n215_})
2'b11 : new_n1167_ = 1'b1;
default : new_n1167_ = 1'b0;
endcase
casez ({u[2], new_n215_})
2'b01 : new_n1168_ = 1'b1;
default : new_n1168_ = 1'b0;
endcase
casez ({y[2], new_n218_})
2'b11 : new_n1169_ = 1'b1;
default : new_n1169_ = 1'b0;
endcase
casez ({new_n98_, new_n220_})
2'b11 : new_n1170_ = 1'b1;
default : new_n1170_ = 1'b0;
endcase
casez ({new_n97_, new_n109_})
2'b10 : new_n1171_ = 1'b1;
default : new_n1171_ = 1'b0;
endcase
casez ({x[2], new_n115_})
2'b11 : new_n1172_ = 1'b1;
default : new_n1172_ = 1'b0;
endcase
casez ({new_n98_, new_n119_})
2'b11 : new_n1173_ = 1'b1;
default : new_n1173_ = 1'b0;
endcase
casez ({y[2], new_n226_})
2'b01 : new_n1174_ = 1'b1;
default : new_n1174_ = 1'b0;
endcase
casez ({new_n97_, new_n119_})
2'b11 : new_n1175_ = 1'b1;
default : new_n1175_ = 1'b0;
endcase
casez ({y[2], new_n123_})
2'b11 : new_n1176_ = 1'b1;
default : new_n1176_ = 1'b0;
endcase
casez ({x[0], new_n126_})
2'b11 : new_n1177_ = 1'b1;
default : new_n1177_ = 1'b0;
endcase
casez ({new_n88_, new_n133_})
2'b11 : new_n1178_ = 1'b1;
default : new_n1178_ = 1'b0;
endcase
casez ({new_n97_, new_n135_})
2'b11 : new_n1179_ = 1'b1;
default : new_n1179_ = 1'b0;
endcase
casez ({u[1], new_n139_})
2'b11 : new_n1180_ = 1'b1;
default : new_n1180_ = 1'b0;
endcase
casez ({u[1], new_n115_})
2'b01 : new_n1181_ = 1'b1;
default : new_n1181_ = 1'b0;
endcase
casez ({new_n89_, new_n116_})
2'b11 : new_n1182_ = 1'b1;
default : new_n1182_ = 1'b0;
endcase
casez ({new_n137_, new_n157_})
2'b00 : new_n1183_ = 1'b1;
default : new_n1183_ = 1'b0;
endcase
casez ({new_n88_, new_n600_, new_n549_, new_n777_})
4'b11?? : new_n1184_ = 1'b1;
4'b??11 : new_n1184_ = 1'b1;
default : new_n1184_ = 1'b0;
endcase
casez ({new_n122_, new_n785_, new_n202_, new_n714_})
4'b11?? : new_n1185_ = 1'b1;
4'b??11 : new_n1185_ = 1'b1;
default : new_n1185_ = 1'b0;
endcase
casez ({new_n448_, new_n501_})
2'b00 : new_n1186_ = 1'b1;
default : new_n1186_ = 1'b0;
endcase
casez ({new_n414_, new_n551_})
2'b00 : new_n1187_ = 1'b1;
default : new_n1187_ = 1'b0;
endcase
casez ({new_n4647_, new_n494_, new_n864_})
3'b1?? : new_n1188_ = 1'b1;
3'b?11 : new_n1188_ = 1'b1;
default : new_n1188_ = 1'b0;
endcase
casez ({x[1], new_n104_, new_n181_})
3'b11? : new_n1189_ = 1'b1;
3'b??0 : new_n1189_ = 1'b1;
default : new_n1189_ = 1'b0;
endcase
casez ({new_n202_, new_n324_, new_n245_, new_n334_})
4'b11?? : new_n1190_ = 1'b1;
4'b??11 : new_n1190_ = 1'b1;
default : new_n1190_ = 1'b0;
endcase
casez ({new_n253_, new_n636_})
2'b00 : new_n1191_ = 1'b1;
default : new_n1191_ = 1'b0;
endcase
casez ({new_n196_, new_n482_, new_n424_, new_n960_})
4'b11?? : new_n1192_ = 1'b1;
4'b??11 : new_n1192_ = 1'b1;
default : new_n1192_ = 1'b0;
endcase
casez ({new_n140_, new_n1003_, new_n307_, new_n367_})
4'b11?? : new_n1193_ = 1'b1;
4'b??11 : new_n1193_ = 1'b1;
default : new_n1193_ = 1'b0;
endcase
casez ({new_n183_, new_n674_})
2'b00 : new_n1194_ = 1'b1;
default : new_n1194_ = 1'b0;
endcase
casez ({new_n225_, new_n380_})
2'b01 : new_n1195_ = 1'b1;
default : new_n1195_ = 1'b0;
endcase
casez ({new_n115_, new_n711_, new_n178_, new_n482_})
4'b11?? : new_n1196_ = 1'b1;
4'b??11 : new_n1196_ = 1'b1;
default : new_n1196_ = 1'b0;
endcase
casez ({new_n340_, new_n377_, new_n378_, new_n441_})
4'b11?? : new_n1197_ = 1'b1;
4'b??11 : new_n1197_ = 1'b1;
default : new_n1197_ = 1'b0;
endcase
casez ({new_n235_, new_n471_, new_n4661_})
3'b11? : new_n1198_ = 1'b1;
3'b??1 : new_n1198_ = 1'b1;
default : new_n1198_ = 1'b0;
endcase
casez ({new_n106_, new_n257_})
2'b11 : new_n1199_ = 1'b1;
default : new_n1199_ = 1'b0;
endcase
casez ({new_n110_, new_n257_})
2'b11 : new_n1200_ = 1'b1;
default : new_n1200_ = 1'b0;
endcase
casez ({new_n85_, new_n271_})
2'b11 : new_n1201_ = 1'b1;
default : new_n1201_ = 1'b0;
endcase
casez ({new_n95_, new_n555_})
2'b11 : new_n1202_ = 1'b1;
default : new_n1202_ = 1'b0;
endcase
casez ({new_n84_, new_n286_})
2'b11 : new_n1203_ = 1'b1;
default : new_n1203_ = 1'b0;
endcase
casez ({new_n88_, new_n294_})
2'b11 : new_n1204_ = 1'b1;
default : new_n1204_ = 1'b0;
endcase
casez ({new_n89_, new_n181_})
2'b10 : new_n1205_ = 1'b1;
default : new_n1205_ = 1'b0;
endcase
casez ({x[0], new_n335_})
2'b11 : new_n1206_ = 1'b1;
default : new_n1206_ = 1'b0;
endcase
casez ({new_n86_, new_n339_})
2'b11 : new_n1207_ = 1'b1;
default : new_n1207_ = 1'b0;
endcase
casez ({new_n186_, new_n194_})
2'b11 : new_n1208_ = 1'b1;
default : new_n1208_ = 1'b0;
endcase
casez ({x[0], new_n352_})
2'b11 : new_n1209_ = 1'b1;
default : new_n1209_ = 1'b0;
endcase
casez ({x[0], new_n352_})
2'b01 : new_n1210_ = 1'b1;
default : new_n1210_ = 1'b0;
endcase
casez ({new_n103_, new_n381_})
2'b11 : new_n1211_ = 1'b1;
default : new_n1211_ = 1'b0;
endcase
casez ({x[0], new_n1024_})
2'b11 : new_n1212_ = 1'b1;
default : new_n1212_ = 1'b0;
endcase
casez ({new_n94_, new_n395_})
2'b11 : new_n1213_ = 1'b1;
default : new_n1213_ = 1'b0;
endcase
casez ({new_n91_, new_n397_})
2'b11 : new_n1214_ = 1'b1;
default : new_n1214_ = 1'b0;
endcase
casez ({u[0], new_n404_})
2'b11 : new_n1215_ = 1'b1;
default : new_n1215_ = 1'b0;
endcase
casez ({new_n88_, new_n407_})
2'b11 : new_n1216_ = 1'b1;
default : new_n1216_ = 1'b0;
endcase
casez ({new_n274_, new_n420_})
2'b11 : new_n1217_ = 1'b1;
default : new_n1217_ = 1'b0;
endcase
casez ({x[0], new_n423_})
2'b11 : new_n1218_ = 1'b1;
default : new_n1218_ = 1'b0;
endcase
casez ({new_n104_, new_n473_})
2'b11 : new_n1219_ = 1'b1;
default : new_n1219_ = 1'b0;
endcase
casez ({new_n106_, new_n250_})
2'b11 : new_n1220_ = 1'b1;
default : new_n1220_ = 1'b0;
endcase
casez ({new_n79_, new_n259_})
2'b11 : new_n1221_ = 1'b1;
default : new_n1221_ = 1'b0;
endcase
casez ({new_n105_, new_n147_})
2'b11 : new_n1222_ = 1'b1;
default : new_n1222_ = 1'b0;
endcase
casez ({new_n89_, new_n282_})
2'b11 : new_n1223_ = 1'b1;
default : new_n1223_ = 1'b0;
endcase
casez ({new_n84_, new_n179_})
2'b11 : new_n1224_ = 1'b1;
default : new_n1224_ = 1'b0;
endcase
casez ({new_n84_, new_n336_})
2'b11 : new_n1225_ = 1'b1;
default : new_n1225_ = 1'b0;
endcase
casez ({new_n179_, new_n198_})
2'b11 : new_n1226_ = 1'b1;
default : new_n1226_ = 1'b0;
endcase
casez ({x[0], new_n366_})
2'b01 : new_n1227_ = 1'b1;
default : new_n1227_ = 1'b0;
endcase
casez ({new_n88_, new_n122_})
2'b11 : new_n1228_ = 1'b1;
default : new_n1228_ = 1'b0;
endcase
casez ({new_n197_, new_n238_})
2'b00 : new_n1229_ = 1'b1;
default : new_n1229_ = 1'b0;
endcase
casez ({new_n208_, new_n775_, new_n238_, new_n462_})
4'b11?? : new_n1230_ = 1'b1;
4'b??11 : new_n1230_ = 1'b1;
default : new_n1230_ = 1'b0;
endcase
casez ({new_n5457_, new_n302_, new_n1148_})
3'b1?? : new_n1231_ = 1'b1;
3'b?01 : new_n1231_ = 1'b1;
default : new_n1231_ = 1'b0;
endcase
casez ({new_n151_, new_n516_, new_n188_, new_n336_})
4'b11?? : new_n1232_ = 1'b1;
4'b??11 : new_n1232_ = 1'b1;
default : new_n1232_ = 1'b0;
endcase
casez ({new_n145_, new_n1182_, new_n151_, new_n696_})
4'b11?? : new_n1233_ = 1'b1;
4'b??11 : new_n1233_ = 1'b1;
default : new_n1233_ = 1'b0;
endcase
casez ({new_n378_, new_n382_, new_n403_, new_n815_})
4'b11?? : new_n1234_ = 1'b1;
4'b??11 : new_n1234_ = 1'b1;
default : new_n1234_ = 1'b0;
endcase
casez ({new_n144_, new_n1216_, new_n224_, new_n464_})
4'b11?? : new_n1235_ = 1'b1;
4'b??11 : new_n1235_ = 1'b1;
default : new_n1235_ = 1'b0;
endcase
casez ({new_n183_, new_n816_, new_n340_, new_n768_})
4'b11?? : new_n1236_ = 1'b1;
4'b??11 : new_n1236_ = 1'b1;
default : new_n1236_ = 1'b0;
endcase
casez ({new_n5454_, new_n350_, new_n462_})
3'b1?? : new_n1237_ = 1'b1;
3'b?11 : new_n1237_ = 1'b1;
default : new_n1237_ = 1'b0;
endcase
casez ({new_n190_, new_n561_, new_n293_, new_n610_})
4'b11?? : new_n1238_ = 1'b1;
4'b??11 : new_n1238_ = 1'b1;
default : new_n1238_ = 1'b0;
endcase
casez ({new_n132_, new_n624_, new_n149_, new_n416_})
4'b11?? : new_n1239_ = 1'b1;
4'b??11 : new_n1239_ = 1'b1;
default : new_n1239_ = 1'b0;
endcase
casez ({new_n176_, new_n464_, new_n5456_})
3'b11? : new_n1240_ = 1'b1;
3'b??1 : new_n1240_ = 1'b1;
default : new_n1240_ = 1'b0;
endcase
casez ({new_n4643_, new_n154_, new_n649_})
3'b1?? : new_n1241_ = 1'b1;
3'b?11 : new_n1241_ = 1'b1;
default : new_n1241_ = 1'b0;
endcase
casez ({new_n80_, new_n269_})
2'b11 : new_n1242_ = 1'b1;
default : new_n1242_ = 1'b0;
endcase
casez ({new_n80_, new_n270_})
2'b11 : new_n1243_ = 1'b1;
default : new_n1243_ = 1'b0;
endcase
casez ({new_n185_, new_n2938_, new_n1184_})
3'b11? : new_n1244_ = 1'b1;
3'b??1 : new_n1244_ = 1'b1;
default : new_n1244_ = 1'b0;
endcase
casez ({new_n95_, new_n1908_, new_n1190_})
3'b11? : new_n1245_ = 1'b1;
3'b??1 : new_n1245_ = 1'b1;
default : new_n1245_ = 1'b0;
endcase
casez ({new_n166_, new_n1923_, new_n1192_})
3'b11? : new_n1246_ = 1'b1;
3'b??1 : new_n1246_ = 1'b1;
default : new_n1246_ = 1'b0;
endcase
casez ({new_n86_, new_n910_, new_n95_, new_n893_})
4'b11?? : new_n1247_ = 1'b1;
4'b??11 : new_n1247_ = 1'b1;
default : new_n1247_ = 1'b0;
endcase
casez ({new_n179_, new_n638_, new_n5927_})
3'b11? : new_n1248_ = 1'b1;
3'b??1 : new_n1248_ = 1'b1;
default : new_n1248_ = 1'b0;
endcase
casez ({new_n115_, new_n693_, new_n293_, new_n704_})
4'b11?? : new_n1249_ = 1'b1;
4'b??11 : new_n1249_ = 1'b1;
default : new_n1249_ = 1'b0;
endcase
casez ({new_n354_, new_n442_})
2'b00 : new_n1250_ = 1'b1;
default : new_n1250_ = 1'b0;
endcase
casez ({new_n179_, new_n2730_, new_n1128_})
3'b11? : new_n1251_ = 1'b1;
3'b??1 : new_n1251_ = 1'b1;
default : new_n1251_ = 1'b0;
endcase
casez ({new_n129_, new_n249_, new_n258_, new_n1033_})
4'b111? : new_n1252_ = 1'b1;
4'b???1 : new_n1252_ = 1'b1;
default : new_n1252_ = 1'b0;
endcase
casez ({u[1], new_n1088_, new_n103_, new_n886_})
4'b01?? : new_n1253_ = 1'b1;
4'b??11 : new_n1253_ = 1'b1;
default : new_n1253_ = 1'b0;
endcase
casez ({y[2], new_n331_})
2'b11 : new_n1254_ = 1'b1;
default : new_n1254_ = 1'b0;
endcase
casez ({new_n373_, new_n2949_, new_n919_})
3'b11? : new_n1255_ = 1'b1;
3'b??1 : new_n1255_ = 1'b1;
default : new_n1255_ = 1'b0;
endcase
casez ({new_n3419_, new_n1255_})
2'b1? : new_n1256_ = 1'b1;
2'b?1 : new_n1256_ = 1'b1;
default : new_n1256_ = 1'b0;
endcase
casez ({u[2], v[1]})
2'b11 : new_n1257_ = 1'b1;
default : new_n1257_ = 1'b0;
endcase
casez ({x[0], u[1]})
2'b01 : new_n1258_ = 1'b1;
default : new_n1258_ = 1'b0;
endcase
casez ({u[2], v[0], new_n2945_})
3'b11? : new_n1259_ = 1'b1;
3'b??1 : new_n1259_ = 1'b1;
default : new_n1259_ = 1'b0;
endcase
casez ({new_n2506_, new_n2519_})
2'b1? : new_n1260_ = 1'b1;
2'b?1 : new_n1260_ = 1'b1;
default : new_n1260_ = 1'b0;
endcase
casez ({new_n284_, new_n305_})
2'b00 : new_n1261_ = 1'b1;
default : new_n1261_ = 1'b0;
endcase
casez ({new_n103_, new_n242_})
2'b00 : new_n1262_ = 1'b1;
default : new_n1262_ = 1'b0;
endcase
casez ({new_n95_, new_n487_})
2'b00 : new_n1263_ = 1'b1;
default : new_n1263_ = 1'b0;
endcase
casez ({new_n86_, new_n88_})
2'b10 : new_n1264_ = 1'b1;
default : new_n1264_ = 1'b0;
endcase
casez ({new_n101_, new_n104_})
2'b11 : new_n1265_ = 1'b1;
default : new_n1265_ = 1'b0;
endcase
casez ({new_n234_, new_n444_})
2'b11 : new_n1266_ = 1'b1;
default : new_n1266_ = 1'b0;
endcase
casez ({x[0], new_n85_})
2'b00 : new_n1267_ = 1'b1;
default : new_n1267_ = 1'b0;
endcase
casez ({y[2], new_n235_, new_n1880_})
3'b11? : new_n1268_ = 1'b1;
3'b??1 : new_n1268_ = 1'b1;
default : new_n1268_ = 1'b0;
endcase
casez ({new_n1639_, new_n2772_})
2'b1? : new_n1269_ = 1'b1;
2'b?1 : new_n1269_ = 1'b1;
default : new_n1269_ = 1'b0;
endcase
casez ({new_n1944_, new_n1629_})
2'b1? : new_n1270_ = 1'b1;
2'b?1 : new_n1270_ = 1'b1;
default : new_n1270_ = 1'b0;
endcase
casez ({new_n2973_, new_n2762_})
2'b1? : new_n1271_ = 1'b1;
2'b?1 : new_n1271_ = 1'b1;
default : new_n1271_ = 1'b0;
endcase
casez ({new_n115_, new_n299_, new_n142_, new_n487_})
4'b11?? : new_n1272_ = 1'b1;
4'b??11 : new_n1272_ = 1'b1;
default : new_n1272_ = 1'b0;
endcase
casez ({v[2], new_n194_, new_n244_, new_n509_})
4'b01?? : new_n1273_ = 1'b1;
4'b??11 : new_n1273_ = 1'b1;
default : new_n1273_ = 1'b0;
endcase
casez ({new_n2602_, new_n254_, new_n531_})
3'b1?? : new_n1274_ = 1'b1;
3'b?11 : new_n1274_ = 1'b1;
default : new_n1274_ = 1'b0;
endcase
casez ({new_n2579_, new_n1588_})
2'b1? : new_n1275_ = 1'b1;
2'b?1 : new_n1275_ = 1'b1;
default : new_n1275_ = 1'b0;
endcase
casez ({new_n205_, new_n532_})
2'b00 : new_n1276_ = 1'b1;
default : new_n1276_ = 1'b0;
endcase
casez ({new_n166_, new_n273_, new_n199_, new_n214_})
4'b11?? : new_n1277_ = 1'b1;
4'b??11 : new_n1277_ = 1'b1;
default : new_n1277_ = 1'b0;
endcase
casez ({new_n3573_, new_n158_, new_n274_})
3'b1?? : new_n1278_ = 1'b1;
3'b?11 : new_n1278_ = 1'b1;
default : new_n1278_ = 1'b0;
endcase
casez ({new_n2693_, new_n3505_})
2'b1? : new_n1279_ = 1'b1;
2'b?1 : new_n1279_ = 1'b1;
default : new_n1279_ = 1'b0;
endcase
casez ({new_n235_, new_n241_, new_n249_, new_n279_})
4'b11?? : new_n1280_ = 1'b1;
4'b??11 : new_n1280_ = 1'b1;
default : new_n1280_ = 1'b0;
endcase
casez ({new_n86_, new_n148_, new_n1947_})
3'b01? : new_n1281_ = 1'b1;
3'b??1 : new_n1281_ = 1'b1;
default : new_n1281_ = 1'b0;
endcase
casez ({new_n91_, new_n124_, new_n190_, new_n284_})
4'b11?? : new_n1282_ = 1'b1;
4'b??11 : new_n1282_ = 1'b1;
default : new_n1282_ = 1'b0;
endcase
casez ({new_n178_, new_n274_, new_n187_, new_n287_})
4'b11?? : new_n1283_ = 1'b1;
4'b??11 : new_n1283_ = 1'b1;
default : new_n1283_ = 1'b0;
endcase
casez ({new_n131_, new_n299_, new_n145_, new_n214_})
4'b11?? : new_n1284_ = 1'b1;
4'b??11 : new_n1284_ = 1'b1;
default : new_n1284_ = 1'b0;
endcase
casez ({new_n1894_, new_n3509_})
2'b1? : new_n1285_ = 1'b1;
2'b?1 : new_n1285_ = 1'b1;
default : new_n1285_ = 1'b0;
endcase
casez ({new_n3481_, new_n155_, new_n166_})
3'b1?? : new_n1286_ = 1'b1;
3'b?11 : new_n1286_ = 1'b1;
default : new_n1286_ = 1'b0;
endcase
casez ({new_n3366_, new_n2572_})
2'b1? : new_n1287_ = 1'b1;
2'b?1 : new_n1287_ = 1'b1;
default : new_n1287_ = 1'b0;
endcase
casez ({new_n3424_, new_n199_, new_n309_})
3'b1?? : new_n1288_ = 1'b1;
3'b?11 : new_n1288_ = 1'b1;
default : new_n1288_ = 1'b0;
endcase
casez ({new_n1625_, new_n84_, new_n598_})
3'b1?? : new_n1289_ = 1'b1;
3'b?11 : new_n1289_ = 1'b1;
default : new_n1289_ = 1'b0;
endcase
casez ({new_n131_, new_n598_, new_n2606_})
3'b11? : new_n1290_ = 1'b1;
3'b??1 : new_n1290_ = 1'b1;
default : new_n1290_ = 1'b0;
endcase
casez ({new_n139_, new_n313_, new_n3334_})
3'b11? : new_n1291_ = 1'b1;
3'b??1 : new_n1291_ = 1'b1;
default : new_n1291_ = 1'b0;
endcase
casez ({new_n3493_, y[2], new_n285_})
3'b1?? : new_n1292_ = 1'b1;
3'b?01 : new_n1292_ = 1'b1;
default : new_n1292_ = 1'b0;
endcase
casez ({new_n194_, new_n315_, new_n2557_})
3'b11? : new_n1293_ = 1'b1;
3'b??1 : new_n1293_ = 1'b1;
default : new_n1293_ = 1'b0;
endcase
casez ({new_n2678_, new_n2512_})
2'b1? : new_n1294_ = 1'b1;
2'b?1 : new_n1294_ = 1'b1;
default : new_n1294_ = 1'b0;
endcase
casez ({new_n3494_, new_n2555_})
2'b1? : new_n1295_ = 1'b1;
2'b?1 : new_n1295_ = 1'b1;
default : new_n1295_ = 1'b0;
endcase
casez ({new_n240_, new_n315_})
2'b00 : new_n1296_ = 1'b1;
default : new_n1296_ = 1'b0;
endcase
casez ({new_n1868_, new_n2718_})
2'b1? : new_n1297_ = 1'b1;
2'b?1 : new_n1297_ = 1'b1;
default : new_n1297_ = 1'b0;
endcase
casez ({new_n1916_, new_n199_, new_n332_})
3'b1?? : new_n1298_ = 1'b1;
3'b?11 : new_n1298_ = 1'b1;
default : new_n1298_ = 1'b0;
endcase
casez ({new_n3413_, new_n191_, new_n332_})
3'b1?? : new_n1299_ = 1'b1;
3'b?11 : new_n1299_ = 1'b1;
default : new_n1299_ = 1'b0;
endcase
casez ({new_n139_, new_n144_, new_n150_, new_n190_})
4'b11?? : new_n1300_ = 1'b1;
4'b??11 : new_n1300_ = 1'b1;
default : new_n1300_ = 1'b0;
endcase
casez ({new_n3490_, new_n1845_})
2'b1? : new_n1301_ = 1'b1;
2'b?1 : new_n1301_ = 1'b1;
default : new_n1301_ = 1'b0;
endcase
casez ({new_n1894_, new_n209_, new_n344_})
3'b1?? : new_n1302_ = 1'b1;
3'b?11 : new_n1302_ = 1'b1;
default : new_n1302_ = 1'b0;
endcase
casez ({new_n183_, new_n199_})
2'b00 : new_n1303_ = 1'b1;
default : new_n1303_ = 1'b0;
endcase
casez ({new_n3480_, new_n2625_})
2'b1? : new_n1304_ = 1'b1;
2'b?1 : new_n1304_ = 1'b1;
default : new_n1304_ = 1'b0;
endcase
casez ({new_n207_, new_n356_})
2'b00 : new_n1305_ = 1'b1;
default : new_n1305_ = 1'b0;
endcase
casez ({new_n140_, new_n356_, new_n3427_})
3'b11? : new_n1306_ = 1'b1;
3'b??1 : new_n1306_ = 1'b1;
default : new_n1306_ = 1'b0;
endcase
casez ({new_n104_, new_n209_, new_n167_, new_n358_})
4'b11?? : new_n1307_ = 1'b1;
4'b??11 : new_n1307_ = 1'b1;
default : new_n1307_ = 1'b0;
endcase
casez ({new_n104_, new_n155_, new_n129_, new_n204_})
4'b11?? : new_n1308_ = 1'b1;
4'b??11 : new_n1308_ = 1'b1;
default : new_n1308_ = 1'b0;
endcase
casez ({new_n3526_, new_n3429_})
2'b1? : new_n1309_ = 1'b1;
2'b?1 : new_n1309_ = 1'b1;
default : new_n1309_ = 1'b0;
endcase
casez ({new_n1830_, new_n3409_})
2'b1? : new_n1310_ = 1'b1;
2'b?1 : new_n1310_ = 1'b1;
default : new_n1310_ = 1'b0;
endcase
casez ({new_n2771_, new_n1851_})
2'b1? : new_n1311_ = 1'b1;
2'b?1 : new_n1311_ = 1'b1;
default : new_n1311_ = 1'b0;
endcase
casez ({new_n144_, new_n194_, new_n1919_})
3'b11? : new_n1312_ = 1'b1;
3'b??1 : new_n1312_ = 1'b1;
default : new_n1312_ = 1'b0;
endcase
casez ({new_n1910_, new_n2634_})
2'b1? : new_n1313_ = 1'b1;
2'b?1 : new_n1313_ = 1'b1;
default : new_n1313_ = 1'b0;
endcase
casez ({new_n1855_, new_n2601_})
2'b1? : new_n1314_ = 1'b1;
2'b?1 : new_n1314_ = 1'b1;
default : new_n1314_ = 1'b0;
endcase
casez ({new_n3423_, new_n98_, new_n123_})
3'b1?? : new_n1315_ = 1'b1;
3'b?01 : new_n1315_ = 1'b1;
default : new_n1315_ = 1'b0;
endcase
casez ({new_n79_, new_n173_, new_n3523_})
3'b11? : new_n1316_ = 1'b1;
3'b??1 : new_n1316_ = 1'b1;
default : new_n1316_ = 1'b0;
endcase
casez ({new_n89_, new_n142_, new_n2734_})
3'b11? : new_n1317_ = 1'b1;
3'b??1 : new_n1317_ = 1'b1;
default : new_n1317_ = 1'b0;
endcase
casez ({new_n2612_, new_n219_, new_n221_})
3'b1?? : new_n1318_ = 1'b1;
3'b?11 : new_n1318_ = 1'b1;
default : new_n1318_ = 1'b0;
endcase
casez ({new_n88_, new_n118_, new_n2662_})
3'b11? : new_n1319_ = 1'b1;
3'b??1 : new_n1319_ = 1'b1;
default : new_n1319_ = 1'b0;
endcase
casez ({new_n137_, new_n411_, new_n209_, new_n226_})
4'b11?? : new_n1320_ = 1'b1;
4'b??11 : new_n1320_ = 1'b1;
default : new_n1320_ = 1'b0;
endcase
casez ({new_n83_, new_n217_, new_n3543_})
3'b01? : new_n1321_ = 1'b1;
3'b??1 : new_n1321_ = 1'b1;
default : new_n1321_ = 1'b0;
endcase
casez ({new_n118_, new_n137_, new_n162_, new_n226_})
4'b11?? : new_n1322_ = 1'b1;
4'b??11 : new_n1322_ = 1'b1;
default : new_n1322_ = 1'b0;
endcase
casez ({new_n79_, new_n120_, new_n91_, new_n115_})
4'b11?? : new_n1323_ = 1'b1;
4'b??11 : new_n1323_ = 1'b1;
default : new_n1323_ = 1'b0;
endcase
casez ({new_n2664_, new_n191_, new_n216_})
3'b1?? : new_n1324_ = 1'b1;
3'b?11 : new_n1324_ = 1'b1;
default : new_n1324_ = 1'b0;
endcase
casez ({new_n3399_, new_n3436_})
2'b1? : new_n1325_ = 1'b1;
2'b?1 : new_n1325_ = 1'b1;
default : new_n1325_ = 1'b0;
endcase
casez ({new_n2764_, new_n2952_})
2'b1? : new_n1326_ = 1'b1;
2'b?1 : new_n1326_ = 1'b1;
default : new_n1326_ = 1'b0;
endcase
casez ({new_n118_, new_n438_, new_n162_, new_n190_})
4'b11?? : new_n1327_ = 1'b1;
4'b??11 : new_n1327_ = 1'b1;
default : new_n1327_ = 1'b0;
endcase
casez ({new_n173_, new_n444_, new_n205_, new_n274_})
4'b11?? : new_n1328_ = 1'b1;
4'b??11 : new_n1328_ = 1'b1;
default : new_n1328_ = 1'b0;
endcase
casez ({new_n2729_, new_n1930_})
2'b1? : new_n1329_ = 1'b1;
2'b?1 : new_n1329_ = 1'b1;
default : new_n1329_ = 1'b0;
endcase
casez ({new_n115_, new_n445_, new_n3476_})
3'b11? : new_n1330_ = 1'b1;
3'b??1 : new_n1330_ = 1'b1;
default : new_n1330_ = 1'b0;
endcase
casez ({new_n1641_, new_n3443_})
2'b1? : new_n1331_ = 1'b1;
2'b?1 : new_n1331_ = 1'b1;
default : new_n1331_ = 1'b0;
endcase
casez ({new_n131_, new_n140_, new_n218_, new_n241_})
4'b11?? : new_n1332_ = 1'b1;
4'b??11 : new_n1332_ = 1'b1;
default : new_n1332_ = 1'b0;
endcase
casez ({new_n137_, new_n241_, new_n3524_})
3'b11? : new_n1333_ = 1'b1;
3'b??1 : new_n1333_ = 1'b1;
default : new_n1333_ = 1'b0;
endcase
casez ({new_n2739_, new_n2672_})
2'b1? : new_n1334_ = 1'b1;
2'b?1 : new_n1334_ = 1'b1;
default : new_n1334_ = 1'b0;
endcase
casez ({new_n84_, new_n2934_, new_n133_})
3'b11? : new_n1335_ = 1'b1;
3'b??1 : new_n1335_ = 1'b1;
default : new_n1335_ = 1'b0;
endcase
casez ({new_n189_, new_n249_, new_n217_, new_n219_})
4'b11?? : new_n1336_ = 1'b1;
4'b??11 : new_n1336_ = 1'b1;
default : new_n1336_ = 1'b0;
endcase
casez ({new_n94_, new_n251_})
2'b11 : new_n1337_ = 1'b1;
default : new_n1337_ = 1'b0;
endcase
casez ({new_n101_, new_n262_})
2'b11 : new_n1338_ = 1'b1;
default : new_n1338_ = 1'b0;
endcase
casez ({new_n145_, new_n153_})
2'b11 : new_n1339_ = 1'b1;
default : new_n1339_ = 1'b0;
endcase
casez ({new_n103_, new_n275_})
2'b11 : new_n1340_ = 1'b1;
default : new_n1340_ = 1'b0;
endcase
casez ({new_n129_, new_n274_})
2'b11 : new_n1341_ = 1'b1;
default : new_n1341_ = 1'b0;
endcase
casez ({new_n150_, new_n278_})
2'b11 : new_n1342_ = 1'b1;
default : new_n1342_ = 1'b0;
endcase
casez ({new_n89_, new_n285_})
2'b11 : new_n1343_ = 1'b1;
default : new_n1343_ = 1'b0;
endcase
casez ({v[2], new_n165_})
2'b11 : new_n1344_ = 1'b1;
default : new_n1344_ = 1'b0;
endcase
casez ({new_n150_, new_n166_})
2'b11 : new_n1345_ = 1'b1;
default : new_n1345_ = 1'b0;
endcase
casez ({new_n131_, new_n170_})
2'b11 : new_n1346_ = 1'b1;
default : new_n1346_ = 1'b0;
endcase
casez ({new_n139_, new_n160_})
2'b11 : new_n1347_ = 1'b1;
default : new_n1347_ = 1'b0;
endcase
casez ({new_n131_, new_n301_})
2'b11 : new_n1348_ = 1'b1;
default : new_n1348_ = 1'b0;
endcase
casez ({new_n140_, new_n177_})
2'b11 : new_n1349_ = 1'b1;
default : new_n1349_ = 1'b0;
endcase
casez ({new_n119_, new_n599_})
2'b11 : new_n1350_ = 1'b1;
default : new_n1350_ = 1'b0;
endcase
casez ({new_n115_, new_n178_})
2'b11 : new_n1351_ = 1'b1;
default : new_n1351_ = 1'b0;
endcase
casez ({new_n177_, new_n317_})
2'b11 : new_n1352_ = 1'b1;
default : new_n1352_ = 1'b0;
endcase
casez ({new_n184_, new_n317_})
2'b11 : new_n1353_ = 1'b1;
default : new_n1353_ = 1'b0;
endcase
casez ({new_n139_, new_n184_})
2'b11 : new_n1354_ = 1'b1;
default : new_n1354_ = 1'b0;
endcase
casez ({new_n142_, new_n337_})
2'b11 : new_n1355_ = 1'b1;
default : new_n1355_ = 1'b0;
endcase
casez ({new_n123_, new_n194_})
2'b11 : new_n1356_ = 1'b1;
default : new_n1356_ = 1'b0;
endcase
casez ({new_n127_, new_n194_})
2'b11 : new_n1357_ = 1'b1;
default : new_n1357_ = 1'b0;
endcase
casez ({new_n127_, new_n343_})
2'b11 : new_n1358_ = 1'b1;
default : new_n1358_ = 1'b0;
endcase
casez ({new_n196_, new_n198_})
2'b11 : new_n1359_ = 1'b1;
default : new_n1359_ = 1'b0;
endcase
casez ({new_n94_, new_n199_})
2'b11 : new_n1360_ = 1'b1;
default : new_n1360_ = 1'b0;
endcase
casez ({new_n131_, new_n200_})
2'b11 : new_n1361_ = 1'b1;
default : new_n1361_ = 1'b0;
endcase
casez ({x[1], new_n200_})
2'b11 : new_n1362_ = 1'b1;
default : new_n1362_ = 1'b0;
endcase
casez ({new_n92_, new_n200_})
2'b01 : new_n1363_ = 1'b1;
default : new_n1363_ = 1'b0;
endcase
casez ({new_n198_, new_n201_})
2'b11 : new_n1364_ = 1'b1;
default : new_n1364_ = 1'b0;
endcase
casez ({new_n210_, new_n369_})
2'b11 : new_n1365_ = 1'b1;
default : new_n1365_ = 1'b0;
endcase
casez ({x[1], new_n208_})
2'b01 : new_n1366_ = 1'b1;
default : new_n1366_ = 1'b0;
endcase
casez ({new_n86_, new_n209_})
2'b11 : new_n1367_ = 1'b1;
default : new_n1367_ = 1'b0;
endcase
casez ({new_n115_, new_n210_})
2'b11 : new_n1368_ = 1'b1;
default : new_n1368_ = 1'b0;
endcase
casez ({new_n194_, new_n210_})
2'b11 : new_n1369_ = 1'b1;
default : new_n1369_ = 1'b0;
endcase
casez ({new_n104_, new_n212_})
2'b11 : new_n1370_ = 1'b1;
default : new_n1370_ = 1'b0;
endcase
casez ({new_n159_, new_n212_})
2'b11 : new_n1371_ = 1'b1;
default : new_n1371_ = 1'b0;
endcase
casez ({new_n137_, new_n216_})
2'b11 : new_n1372_ = 1'b1;
default : new_n1372_ = 1'b0;
endcase
casez ({y[2], new_n218_})
2'b01 : new_n1373_ = 1'b1;
default : new_n1373_ = 1'b0;
endcase
casez ({new_n219_, new_n220_})
2'b11 : new_n1374_ = 1'b1;
default : new_n1374_ = 1'b0;
endcase
casez ({new_n215_, new_n228_})
2'b11 : new_n1375_ = 1'b1;
default : new_n1375_ = 1'b0;
endcase
casez ({new_n191_, new_n228_})
2'b11 : new_n1376_ = 1'b1;
default : new_n1376_ = 1'b0;
endcase
casez ({new_n94_, new_n237_})
2'b11 : new_n1377_ = 1'b1;
default : new_n1377_ = 1'b0;
endcase
casez ({new_n94_, new_n120_})
2'b11 : new_n1378_ = 1'b1;
default : new_n1378_ = 1'b0;
endcase
casez ({new_n94_, new_n128_})
2'b11 : new_n1379_ = 1'b1;
default : new_n1379_ = 1'b0;
endcase
casez ({new_n127_, new_n238_})
2'b11 : new_n1380_ = 1'b1;
default : new_n1380_ = 1'b0;
endcase
casez ({new_n154_, new_n239_})
2'b11 : new_n1381_ = 1'b1;
default : new_n1381_ = 1'b0;
endcase
casez ({new_n82_, new_n130_})
2'b01 : new_n1382_ = 1'b1;
default : new_n1382_ = 1'b0;
endcase
casez ({new_n115_, new_n242_})
2'b11 : new_n1383_ = 1'b1;
default : new_n1383_ = 1'b0;
endcase
casez ({new_n151_, new_n243_})
2'b11 : new_n1384_ = 1'b1;
default : new_n1384_ = 1'b0;
endcase
casez ({new_n84_, new_n143_})
2'b11 : new_n1385_ = 1'b1;
default : new_n1385_ = 1'b0;
endcase
casez ({x[0], new_n145_})
2'b01 : new_n1386_ = 1'b1;
default : new_n1386_ = 1'b0;
endcase
casez ({y[2], new_n145_})
2'b01 : new_n1387_ = 1'b1;
default : new_n1387_ = 1'b0;
endcase
casez ({x[2], new_n150_})
2'b01 : new_n1388_ = 1'b1;
default : new_n1388_ = 1'b0;
endcase
casez ({new_n84_, new_n152_})
2'b11 : new_n1389_ = 1'b1;
default : new_n1389_ = 1'b0;
endcase
casez ({new_n98_, new_n152_})
2'b11 : new_n1390_ = 1'b1;
default : new_n1390_ = 1'b0;
endcase
casez ({new_n95_, new_n148_})
2'b11 : new_n1391_ = 1'b1;
default : new_n1391_ = 1'b0;
endcase
casez ({x[2], new_n169_})
2'b01 : new_n1392_ = 1'b1;
default : new_n1392_ = 1'b0;
endcase
casez ({new_n92_, new_n170_})
2'b11 : new_n1393_ = 1'b1;
default : new_n1393_ = 1'b0;
endcase
casez ({y[2], new_n173_})
2'b11 : new_n1394_ = 1'b1;
default : new_n1394_ = 1'b0;
endcase
casez ({u[2], new_n178_})
2'b01 : new_n1395_ = 1'b1;
default : new_n1395_ = 1'b0;
endcase
casez ({new_n93_, new_n177_})
2'b11 : new_n1396_ = 1'b1;
default : new_n1396_ = 1'b0;
endcase
casez ({u[2], new_n178_})
2'b11 : new_n1397_ = 1'b1;
default : new_n1397_ = 1'b0;
endcase
casez ({new_n92_, new_n187_})
2'b11 : new_n1398_ = 1'b1;
default : new_n1398_ = 1'b0;
endcase
casez ({y[2], new_n189_})
2'b11 : new_n1399_ = 1'b1;
default : new_n1399_ = 1'b0;
endcase
casez ({v[1], new_n190_})
2'b01 : new_n1400_ = 1'b1;
default : new_n1400_ = 1'b0;
endcase
casez ({new_n92_, new_n201_})
2'b01 : new_n1401_ = 1'b1;
default : new_n1401_ = 1'b0;
endcase
casez ({x[2], new_n118_})
2'b01 : new_n1402_ = 1'b1;
default : new_n1402_ = 1'b0;
endcase
casez ({y[2], new_n226_})
2'b11 : new_n1403_ = 1'b1;
default : new_n1403_ = 1'b0;
endcase
casez ({new_n371_, new_n768_})
2'b00 : new_n1404_ = 1'b1;
default : new_n1404_ = 1'b0;
endcase
casez ({new_n129_, new_n253_})
2'b00 : new_n1405_ = 1'b1;
default : new_n1405_ = 1'b0;
endcase
casez ({new_n86_, new_n495_, new_n4668_})
3'b11? : new_n1406_ = 1'b1;
3'b??1 : new_n1406_ = 1'b1;
default : new_n1406_ = 1'b0;
endcase
casez ({new_n2811_, new_n2694_})
2'b1? : new_n1407_ = 1'b1;
2'b?1 : new_n1407_ = 1'b1;
default : new_n1407_ = 1'b0;
endcase
casez ({new_n4641_, new_n157_, new_n211_})
3'b1?? : new_n1408_ = 1'b1;
3'b?11 : new_n1408_ = 1'b1;
default : new_n1408_ = 1'b0;
endcase
casez ({new_n280_, new_n787_})
2'b00 : new_n1409_ = 1'b1;
default : new_n1409_ = 1'b0;
endcase
casez ({new_n93_, new_n502_, new_n144_, new_n356_})
4'b11?? : new_n1410_ = 1'b1;
4'b??11 : new_n1410_ = 1'b1;
default : new_n1410_ = 1'b0;
endcase
casez ({new_n2846_, new_n157_, new_n264_})
3'b1?? : new_n1411_ = 1'b1;
3'b?11 : new_n1411_ = 1'b1;
default : new_n1411_ = 1'b0;
endcase
casez ({new_n414_, new_n797_})
2'b00 : new_n1412_ = 1'b1;
default : new_n1412_ = 1'b0;
endcase
casez ({new_n405_, new_n800_})
2'b00 : new_n1413_ = 1'b1;
default : new_n1413_ = 1'b0;
endcase
casez ({new_n2111_, new_n2660_})
2'b1? : new_n1414_ = 1'b1;
2'b?1 : new_n1414_ = 1'b1;
default : new_n1414_ = 1'b0;
endcase
casez ({new_n2113_, new_n3367_})
2'b1? : new_n1415_ = 1'b1;
2'b?1 : new_n1415_ = 1'b1;
default : new_n1415_ = 1'b0;
endcase
casez ({new_n1718_, new_n1719_})
2'b1? : new_n1416_ = 1'b1;
2'b?1 : new_n1416_ = 1'b1;
default : new_n1416_ = 1'b0;
endcase
casez ({new_n2817_, new_n2686_})
2'b1? : new_n1417_ = 1'b1;
2'b?1 : new_n1417_ = 1'b1;
default : new_n1417_ = 1'b0;
endcase
casez ({new_n93_, new_n280_, new_n1919_})
3'b11? : new_n1418_ = 1'b1;
3'b??1 : new_n1418_ = 1'b1;
default : new_n1418_ = 1'b0;
endcase
casez ({new_n96_, new_n282_, new_n131_, new_n192_})
4'b11?? : new_n1419_ = 1'b1;
4'b??11 : new_n1419_ = 1'b1;
default : new_n1419_ = 1'b0;
endcase
casez ({new_n104_, new_n553_, new_n380_, new_n527_})
4'b01?? : new_n1420_ = 1'b1;
4'b??01 : new_n1420_ = 1'b1;
default : new_n1420_ = 1'b0;
endcase
casez ({new_n115_, new_n555_, new_n131_, new_n483_})
4'b11?? : new_n1421_ = 1'b1;
4'b??11 : new_n1421_ = 1'b1;
default : new_n1421_ = 1'b0;
endcase
casez ({new_n101_, new_n295_, new_n118_, new_n215_})
4'b11?? : new_n1422_ = 1'b1;
4'b??11 : new_n1422_ = 1'b1;
default : new_n1422_ = 1'b0;
endcase
casez ({new_n268_, new_n872_})
2'b00 : new_n1423_ = 1'b1;
default : new_n1423_ = 1'b0;
endcase
casez ({new_n104_, new_n1344_, new_n144_, new_n159_})
4'b11?? : new_n1424_ = 1'b1;
4'b??11 : new_n1424_ = 1'b1;
default : new_n1424_ = 1'b0;
endcase
casez ({new_n2822_, new_n153_, new_n293_})
3'b1?? : new_n1425_ = 1'b1;
3'b?11 : new_n1425_ = 1'b1;
default : new_n1425_ = 1'b0;
endcase
casez ({y[2], new_n606_, new_n4655_})
3'b01? : new_n1426_ = 1'b1;
3'b??1 : new_n1426_ = 1'b1;
default : new_n1426_ = 1'b0;
endcase
casez ({new_n4605_, new_n3466_})
2'b1? : new_n1427_ = 1'b1;
2'b?1 : new_n1427_ = 1'b1;
default : new_n1427_ = 1'b0;
endcase
casez ({new_n2603_, new_n243_, new_n359_})
3'b1?? : new_n1428_ = 1'b1;
3'b?10 : new_n1428_ = 1'b1;
default : new_n1428_ = 1'b0;
endcase
casez ({new_n3435_, new_n672_})
2'b1? : new_n1429_ = 1'b1;
2'b?1 : new_n1429_ = 1'b1;
default : new_n1429_ = 1'b0;
endcase
casez ({v[1], new_n2933_, new_n673_})
3'b01? : new_n1430_ = 1'b1;
3'b??1 : new_n1430_ = 1'b1;
default : new_n1430_ = 1'b0;
endcase
casez ({new_n2138_, new_n144_, new_n281_})
3'b1?? : new_n1431_ = 1'b1;
3'b?11 : new_n1431_ = 1'b1;
default : new_n1431_ = 1'b0;
endcase
casez ({new_n4664_, new_n115_, new_n229_})
3'b1?? : new_n1432_ = 1'b1;
3'b?11 : new_n1432_ = 1'b1;
default : new_n1432_ = 1'b0;
endcase
casez ({new_n577_, new_n1011_})
2'b00 : new_n1433_ = 1'b1;
default : new_n1433_ = 1'b0;
endcase
casez ({new_n4656_, new_n2641_})
2'b1? : new_n1434_ = 1'b1;
2'b?1 : new_n1434_ = 1'b1;
default : new_n1434_ = 1'b0;
endcase
casez ({new_n4656_, new_n131_, new_n229_})
3'b1?? : new_n1435_ = 1'b1;
3'b?11 : new_n1435_ = 1'b1;
default : new_n1435_ = 1'b0;
endcase
casez ({new_n2831_, new_n2694_})
2'b1? : new_n1436_ = 1'b1;
2'b?1 : new_n1436_ = 1'b1;
default : new_n1436_ = 1'b0;
endcase
casez ({v[0], new_n680_, new_n3372_})
3'b01? : new_n1437_ = 1'b1;
3'b??1 : new_n1437_ = 1'b1;
default : new_n1437_ = 1'b0;
endcase
casez ({new_n780_, new_n1018_})
2'b00 : new_n1438_ = 1'b1;
default : new_n1438_ = 1'b0;
endcase
casez ({new_n94_, new_n212_, new_n175_, new_n216_})
4'b11?? : new_n1439_ = 1'b1;
4'b??11 : new_n1439_ = 1'b1;
default : new_n1439_ = 1'b0;
endcase
casez ({new_n4658_, new_n1725_})
2'b1? : new_n1440_ = 1'b1;
2'b?1 : new_n1440_ = 1'b1;
default : new_n1440_ = 1'b0;
endcase
casez ({new_n3384_, new_n1733_})
2'b1? : new_n1441_ = 1'b1;
2'b?1 : new_n1441_ = 1'b1;
default : new_n1441_ = 1'b0;
endcase
casez ({new_n118_, new_n308_, new_n4620_})
3'b11? : new_n1442_ = 1'b1;
3'b??1 : new_n1442_ = 1'b1;
default : new_n1442_ = 1'b0;
endcase
casez ({new_n81_, new_n398_, new_n261_, new_n332_})
4'b11?? : new_n1443_ = 1'b1;
4'b??11 : new_n1443_ = 1'b1;
default : new_n1443_ = 1'b0;
endcase
casez ({new_n118_, new_n397_, new_n243_, new_n408_})
4'b11?? : new_n1444_ = 1'b1;
4'b??11 : new_n1444_ = 1'b1;
default : new_n1444_ = 1'b0;
endcase
casez ({new_n115_, new_n397_, new_n211_, new_n408_})
4'b11?? : new_n1445_ = 1'b1;
4'b??11 : new_n1445_ = 1'b1;
default : new_n1445_ = 1'b0;
endcase
casez ({new_n3471_, new_n83_, new_n707_})
3'b1?? : new_n1446_ = 1'b1;
3'b?10 : new_n1446_ = 1'b1;
default : new_n1446_ = 1'b0;
endcase
casez ({new_n448_, new_n714_})
2'b00 : new_n1447_ = 1'b1;
default : new_n1447_ = 1'b0;
endcase
casez ({new_n1742_, new_n169_, new_n189_})
3'b1?? : new_n1448_ = 1'b1;
3'b?11 : new_n1448_ = 1'b1;
default : new_n1448_ = 1'b0;
endcase
casez ({new_n450_, new_n717_})
2'b00 : new_n1449_ = 1'b1;
default : new_n1449_ = 1'b0;
endcase
casez ({new_n96_, new_n340_, new_n101_, new_n429_})
4'b11?? : new_n1450_ = 1'b1;
4'b??11 : new_n1450_ = 1'b1;
default : new_n1450_ = 1'b0;
endcase
casez ({new_n120_, new_n177_, new_n204_, new_n442_})
4'b11?? : new_n1451_ = 1'b1;
4'b??11 : new_n1451_ = 1'b1;
default : new_n1451_ = 1'b0;
endcase
casez ({y[2], new_n396_, new_n161_, new_n444_})
4'b01?? : new_n1452_ = 1'b1;
4'b??11 : new_n1452_ = 1'b1;
default : new_n1452_ = 1'b0;
endcase
casez ({y[2], new_n236_, new_n1930_})
3'b01? : new_n1453_ = 1'b1;
3'b??1 : new_n1453_ = 1'b1;
default : new_n1453_ = 1'b0;
endcase
casez ({new_n93_, new_n158_, new_n448_})
3'b01? : new_n1454_ = 1'b1;
3'b??1 : new_n1454_ = 1'b1;
default : new_n1454_ = 1'b0;
endcase
casez ({new_n325_, new_n743_})
2'b00 : new_n1455_ = 1'b1;
default : new_n1455_ = 1'b0;
endcase
casez ({new_n97_, new_n1126_, new_n3428_})
3'b11? : new_n1456_ = 1'b1;
3'b??1 : new_n1456_ = 1'b1;
default : new_n1456_ = 1'b0;
endcase
casez ({new_n112_, new_n260_})
2'b11 : new_n1457_ = 1'b1;
default : new_n1457_ = 1'b0;
endcase
casez ({v[0], new_n526_})
2'b11 : new_n1458_ = 1'b1;
default : new_n1458_ = 1'b0;
endcase
casez ({new_n92_, new_n272_})
2'b11 : new_n1459_ = 1'b1;
default : new_n1459_ = 1'b0;
endcase
casez ({x[0], new_n282_})
2'b01 : new_n1460_ = 1'b1;
default : new_n1460_ = 1'b0;
endcase
casez ({x[0], new_n282_})
2'b11 : new_n1461_ = 1'b1;
default : new_n1461_ = 1'b0;
endcase
casez ({y[2], new_n292_})
2'b01 : new_n1462_ = 1'b1;
default : new_n1462_ = 1'b0;
endcase
casez ({u[0], new_n294_})
2'b11 : new_n1463_ = 1'b1;
default : new_n1463_ = 1'b0;
endcase
casez ({new_n106_, new_n169_})
2'b11 : new_n1464_ = 1'b1;
default : new_n1464_ = 1'b0;
endcase
casez ({new_n89_, new_n581_})
2'b11 : new_n1465_ = 1'b1;
default : new_n1465_ = 1'b0;
endcase
casez ({x[0], new_n310_})
2'b01 : new_n1466_ = 1'b1;
default : new_n1466_ = 1'b0;
endcase
casez ({new_n88_, new_n310_})
2'b11 : new_n1467_ = 1'b1;
default : new_n1467_ = 1'b0;
endcase
casez ({y[2], new_n324_})
2'b11 : new_n1468_ = 1'b1;
default : new_n1468_ = 1'b0;
endcase
casez ({new_n79_, new_n325_})
2'b11 : new_n1469_ = 1'b1;
default : new_n1469_ = 1'b0;
endcase
casez ({new_n77_, new_n329_})
2'b01 : new_n1470_ = 1'b1;
default : new_n1470_ = 1'b0;
endcase
casez ({v[2], new_n329_})
2'b01 : new_n1471_ = 1'b1;
default : new_n1471_ = 1'b0;
endcase
casez ({new_n95_, new_n329_})
2'b11 : new_n1472_ = 1'b1;
default : new_n1472_ = 1'b0;
endcase
casez ({new_n86_, new_n330_})
2'b11 : new_n1473_ = 1'b1;
default : new_n1473_ = 1'b0;
endcase
casez ({u[0], new_n352_})
2'b11 : new_n1474_ = 1'b1;
default : new_n1474_ = 1'b0;
endcase
casez ({new_n96_, new_n352_})
2'b11 : new_n1475_ = 1'b1;
default : new_n1475_ = 1'b0;
endcase
casez ({u[0], new_n352_})
2'b01 : new_n1476_ = 1'b1;
default : new_n1476_ = 1'b0;
endcase
casez ({new_n92_, new_n202_})
2'b11 : new_n1477_ = 1'b1;
default : new_n1477_ = 1'b0;
endcase
casez ({new_n89_, new_n366_})
2'b11 : new_n1478_ = 1'b1;
default : new_n1478_ = 1'b0;
endcase
casez ({new_n89_, new_n382_})
2'b11 : new_n1479_ = 1'b1;
default : new_n1479_ = 1'b0;
endcase
casez ({new_n96_, new_n383_})
2'b11 : new_n1480_ = 1'b1;
default : new_n1480_ = 1'b0;
endcase
casez ({new_n170_, new_n388_})
2'b11 : new_n1481_ = 1'b1;
default : new_n1481_ = 1'b0;
endcase
casez ({new_n178_, new_n388_})
2'b11 : new_n1482_ = 1'b1;
default : new_n1482_ = 1'b0;
endcase
casez ({new_n103_, new_n389_})
2'b11 : new_n1483_ = 1'b1;
default : new_n1483_ = 1'b0;
endcase
casez ({x[0], new_n407_})
2'b11 : new_n1484_ = 1'b1;
default : new_n1484_ = 1'b0;
endcase
casez ({new_n91_, new_n408_})
2'b11 : new_n1485_ = 1'b1;
default : new_n1485_ = 1'b0;
endcase
casez ({v[1], new_n422_})
2'b01 : new_n1486_ = 1'b1;
default : new_n1486_ = 1'b0;
endcase
casez ({x[0], new_n429_})
2'b11 : new_n1487_ = 1'b1;
default : new_n1487_ = 1'b0;
endcase
casez ({u[0], new_n429_})
2'b11 : new_n1488_ = 1'b1;
default : new_n1488_ = 1'b0;
endcase
casez ({new_n94_, new_n449_})
2'b11 : new_n1489_ = 1'b1;
default : new_n1489_ = 1'b0;
endcase
casez ({new_n89_, new_n451_})
2'b11 : new_n1490_ = 1'b1;
default : new_n1490_ = 1'b0;
endcase
casez ({new_n79_, new_n458_})
2'b11 : new_n1491_ = 1'b1;
default : new_n1491_ = 1'b0;
endcase
casez ({new_n96_, new_n459_})
2'b11 : new_n1492_ = 1'b1;
default : new_n1492_ = 1'b0;
endcase
casez ({new_n168_, new_n1492_, new_n170_, new_n548_})
4'b11?? : new_n1493_ = 1'b1;
4'b??11 : new_n1493_ = 1'b1;
default : new_n1493_ = 1'b0;
endcase
casez ({new_n102_, new_n136_})
2'b11 : new_n1494_ = 1'b1;
default : new_n1494_ = 1'b0;
endcase
casez ({y[2], new_n472_})
2'b11 : new_n1495_ = 1'b1;
default : new_n1495_ = 1'b0;
endcase
casez ({new_n89_, new_n157_})
2'b11 : new_n1496_ = 1'b1;
default : new_n1496_ = 1'b0;
endcase
casez ({new_n88_, new_n282_})
2'b11 : new_n1497_ = 1'b1;
default : new_n1497_ = 1'b0;
endcase
casez ({new_n84_, new_n268_})
2'b11 : new_n1498_ = 1'b1;
default : new_n1498_ = 1'b0;
endcase
casez ({new_n79_, new_n303_})
2'b11 : new_n1499_ = 1'b1;
default : new_n1499_ = 1'b0;
endcase
casez ({u[0], new_n335_})
2'b01 : new_n1500_ = 1'b1;
default : new_n1500_ = 1'b0;
endcase
casez ({new_n101_, new_n383_})
2'b11 : new_n1501_ = 1'b1;
default : new_n1501_ = 1'b0;
endcase
casez ({new_n96_, new_n390_})
2'b11 : new_n1502_ = 1'b1;
default : new_n1502_ = 1'b0;
endcase
casez ({new_n83_, new_n113_})
2'b11 : new_n1503_ = 1'b1;
default : new_n1503_ = 1'b0;
endcase
casez ({new_n85_, new_n114_})
2'b11 : new_n1504_ = 1'b1;
default : new_n1504_ = 1'b0;
endcase
casez ({x[0], new_n459_})
2'b01 : new_n1505_ = 1'b1;
default : new_n1505_ = 1'b0;
endcase
casez ({new_n195_, new_n197_})
2'b00 : new_n1506_ = 1'b1;
default : new_n1506_ = 1'b0;
endcase
casez ({new_n83_, new_n149_, new_n3517_})
3'b11? : new_n1507_ = 1'b1;
3'b??1 : new_n1507_ = 1'b1;
default : new_n1507_ = 1'b0;
endcase
casez ({new_n164_, new_n444_, new_n168_, new_n411_})
4'b11?? : new_n1508_ = 1'b1;
4'b??11 : new_n1508_ = 1'b1;
default : new_n1508_ = 1'b0;
endcase
casez ({new_n96_, new_n1199_, new_n274_, new_n389_})
4'b01?? : new_n1509_ = 1'b1;
4'b??11 : new_n1509_ = 1'b1;
default : new_n1509_ = 1'b0;
endcase
casez ({new_n5453_, new_n129_, new_n194_})
3'b1?? : new_n1510_ = 1'b1;
3'b?11 : new_n1510_ = 1'b1;
default : new_n1510_ = 1'b0;
endcase
casez ({new_n3444_, new_n825_})
2'b1? : new_n1511_ = 1'b1;
2'b?1 : new_n1511_ = 1'b1;
default : new_n1511_ = 1'b0;
endcase
casez ({new_n97_, new_n283_, new_n182_, new_n287_})
4'b11?? : new_n1512_ = 1'b1;
4'b??11 : new_n1512_ = 1'b1;
default : new_n1512_ = 1'b0;
endcase
casez ({new_n512_, new_n567_})
2'b00 : new_n1513_ = 1'b1;
default : new_n1513_ = 1'b0;
endcase
casez ({new_n182_, new_n571_})
2'b00 : new_n1514_ = 1'b1;
default : new_n1514_ = 1'b0;
endcase
casez ({new_n870_, new_n900_})
2'b00 : new_n1515_ = 1'b1;
default : new_n1515_ = 1'b0;
endcase
casez ({new_n696_, new_n903_})
2'b00 : new_n1516_ = 1'b1;
default : new_n1516_ = 1'b0;
endcase
casez ({u[2], new_n312_, new_n80_, new_n637_})
4'b01?? : new_n1517_ = 1'b1;
4'b??01 : new_n1517_ = 1'b1;
default : new_n1517_ = 1'b0;
endcase
casez ({new_n89_, new_n164_, new_n121_, new_n344_})
4'b11?? : new_n1518_ = 1'b1;
4'b??11 : new_n1518_ = 1'b1;
default : new_n1518_ = 1'b0;
endcase
casez ({y[2], new_n734_, new_n153_, new_n656_})
4'b11?? : new_n1519_ = 1'b1;
4'b??11 : new_n1519_ = 1'b1;
default : new_n1519_ = 1'b0;
endcase
casez ({new_n384_, new_n463_})
2'b00 : new_n1520_ = 1'b1;
default : new_n1520_ = 1'b0;
endcase
casez ({u[0], new_n168_, new_n3557_})
3'b01? : new_n1521_ = 1'b1;
3'b??1 : new_n1521_ = 1'b1;
default : new_n1521_ = 1'b0;
endcase
casez ({new_n164_, new_n249_, new_n168_, new_n241_})
4'b11?? : new_n1522_ = 1'b1;
4'b??11 : new_n1522_ = 1'b1;
default : new_n1522_ = 1'b0;
endcase
casez ({new_n97_, new_n277_})
2'b11 : new_n1523_ = 1'b1;
default : new_n1523_ = 1'b0;
endcase
casez ({v[1], new_n283_})
2'b11 : new_n1524_ = 1'b1;
default : new_n1524_ = 1'b0;
endcase
casez ({y[2], new_n168_})
2'b01 : new_n1525_ = 1'b1;
default : new_n1525_ = 1'b0;
endcase
casez ({new_n373_, new_n401_})
2'b11 : new_n1526_ = 1'b1;
default : new_n1526_ = 1'b0;
endcase
casez ({new_n5926_, new_n248_, new_n775_})
3'b1?? : new_n1527_ = 1'b1;
3'b?11 : new_n1527_ = 1'b1;
default : new_n1527_ = 1'b0;
endcase
casez ({new_n592_, new_n870_})
2'b00 : new_n1528_ = 1'b1;
default : new_n1528_ = 1'b0;
endcase
casez ({new_n585_, new_n889_})
2'b00 : new_n1529_ = 1'b1;
default : new_n1529_ = 1'b0;
endcase
casez ({y[2], new_n608_, new_n1905_})
3'b01? : new_n1530_ = 1'b1;
3'b??1 : new_n1530_ = 1'b1;
default : new_n1530_ = 1'b0;
endcase
casez ({new_n97_, new_n1882_, new_n1426_})
3'b11? : new_n1531_ = 1'b1;
3'b??1 : new_n1531_ = 1'b1;
default : new_n1531_ = 1'b0;
endcase
casez ({new_n193_, new_n597_, new_n304_, new_n1506_})
4'b11?? : new_n1532_ = 1'b1;
4'b??00 : new_n1532_ = 1'b1;
default : new_n1532_ = 1'b0;
endcase
casez ({new_n440_, new_n804_})
2'b00 : new_n1533_ = 1'b1;
default : new_n1533_ = 1'b0;
endcase
casez ({new_n415_, new_n977_})
2'b00 : new_n1534_ = 1'b1;
default : new_n1534_ = 1'b0;
endcase
casez ({new_n563_, new_n703_})
2'b00 : new_n1535_ = 1'b1;
default : new_n1535_ = 1'b0;
endcase
casez ({new_n280_, new_n704_})
2'b00 : new_n1536_ = 1'b1;
default : new_n1536_ = 1'b0;
endcase
casez ({new_n86_, new_n117_, new_n196_, new_n235_})
4'b11?? : new_n1537_ = 1'b1;
4'b??11 : new_n1537_ = 1'b1;
default : new_n1537_ = 1'b0;
endcase
casez ({u[2], new_n298_, new_n113_, new_n198_})
4'b11?? : new_n1538_ = 1'b1;
4'b??11 : new_n1538_ = 1'b1;
default : new_n1538_ = 1'b0;
endcase
casez ({v[0], v[2]})
2'b11 : new_n1539_ = 1'b1;
default : new_n1539_ = 1'b0;
endcase
casez ({new_n86_, new_n284_})
2'b00 : new_n1540_ = 1'b1;
default : new_n1540_ = 1'b0;
endcase
casez ({new_n89_, new_n224_})
2'b00 : new_n1541_ = 1'b1;
default : new_n1541_ = 1'b0;
endcase
casez ({new_n93_, new_n103_})
2'b11 : new_n1542_ = 1'b1;
default : new_n1542_ = 1'b0;
endcase
casez ({new_n93_, new_n104_})
2'b11 : new_n1543_ = 1'b1;
default : new_n1543_ = 1'b0;
endcase
casez ({new_n86_, new_n101_})
2'b01 : new_n1544_ = 1'b1;
default : new_n1544_ = 1'b0;
endcase
casez ({u[0], new_n103_})
2'b10 : new_n1545_ = 1'b1;
default : new_n1545_ = 1'b0;
endcase
casez ({new_n80_, new_n86_})
2'b11 : new_n1546_ = 1'b1;
default : new_n1546_ = 1'b0;
endcase
casez ({new_n144_, new_n155_})
2'b00 : new_n1547_ = 1'b1;
default : new_n1547_ = 1'b0;
endcase
casez ({new_n346_, new_n564_})
2'b01 : new_n1548_ = 1'b1;
default : new_n1548_ = 1'b0;
endcase
casez ({new_n248_, new_n293_})
2'b00 : new_n1549_ = 1'b1;
default : new_n1549_ = 1'b0;
endcase
casez ({new_n174_, new_n926_})
2'b00 : new_n1550_ = 1'b1;
default : new_n1550_ = 1'b0;
endcase
casez ({new_n2511_, new_n342_})
2'b1? : new_n1551_ = 1'b1;
2'b?1 : new_n1551_ = 1'b1;
default : new_n1551_ = 1'b0;
endcase
casez ({new_n254_, new_n344_})
2'b00 : new_n1552_ = 1'b1;
default : new_n1552_ = 1'b0;
endcase
casez ({new_n3507_, new_n1098_})
2'b1? : new_n1553_ = 1'b1;
2'b?1 : new_n1553_ = 1'b1;
default : new_n1553_ = 1'b0;
endcase
casez ({new_n212_, new_n250_})
2'b00 : new_n1554_ = 1'b1;
default : new_n1554_ = 1'b0;
endcase
casez ({new_n129_, new_n148_})
2'b11 : new_n1555_ = 1'b1;
default : new_n1555_ = 1'b0;
endcase
casez ({new_n137_, new_n153_})
2'b11 : new_n1556_ = 1'b1;
default : new_n1556_ = 1'b0;
endcase
casez ({u[1], new_n275_})
2'b11 : new_n1557_ = 1'b1;
default : new_n1557_ = 1'b0;
endcase
casez ({new_n131_, new_n281_})
2'b11 : new_n1558_ = 1'b1;
default : new_n1558_ = 1'b0;
endcase
casez ({new_n144_, new_n178_})
2'b11 : new_n1559_ = 1'b1;
default : new_n1559_ = 1'b0;
endcase
casez ({new_n208_, new_n316_})
2'b11 : new_n1560_ = 1'b1;
default : new_n1560_ = 1'b0;
endcase
casez ({new_n145_, new_n332_})
2'b11 : new_n1561_ = 1'b1;
default : new_n1561_ = 1'b0;
endcase
casez ({new_n140_, new_n332_})
2'b11 : new_n1562_ = 1'b1;
default : new_n1562_ = 1'b0;
endcase
casez ({new_n158_, new_n338_})
2'b11 : new_n1563_ = 1'b1;
default : new_n1563_ = 1'b0;
endcase
casez ({new_n161_, new_n338_})
2'b11 : new_n1564_ = 1'b1;
default : new_n1564_ = 1'b0;
endcase
casez ({new_n176_, new_n338_})
2'b11 : new_n1565_ = 1'b1;
default : new_n1565_ = 1'b0;
endcase
casez ({new_n92_, new_n196_})
2'b01 : new_n1566_ = 1'b1;
default : new_n1566_ = 1'b0;
endcase
casez ({new_n93_, new_n201_})
2'b01 : new_n1567_ = 1'b1;
default : new_n1567_ = 1'b0;
endcase
casez ({new_n87_, new_n204_})
2'b11 : new_n1568_ = 1'b1;
default : new_n1568_ = 1'b0;
endcase
casez ({new_n155_, new_n363_})
2'b11 : new_n1569_ = 1'b1;
default : new_n1569_ = 1'b0;
endcase
casez ({new_n79_, new_n206_})
2'b01 : new_n1570_ = 1'b1;
default : new_n1570_ = 1'b0;
endcase
casez ({new_n212_, new_n220_})
2'b11 : new_n1571_ = 1'b1;
default : new_n1571_ = 1'b0;
endcase
casez ({new_n115_, new_n223_})
2'b11 : new_n1572_ = 1'b1;
default : new_n1572_ = 1'b0;
endcase
casez ({new_n166_, new_n417_})
2'b11 : new_n1573_ = 1'b1;
default : new_n1573_ = 1'b0;
endcase
casez ({new_n154_, new_n228_})
2'b11 : new_n1574_ = 1'b1;
default : new_n1574_ = 1'b0;
endcase
casez ({v[2], new_n120_})
2'b01 : new_n1575_ = 1'b1;
default : new_n1575_ = 1'b0;
endcase
casez ({new_n170_, new_n432_})
2'b11 : new_n1576_ = 1'b1;
default : new_n1576_ = 1'b0;
endcase
casez ({new_n84_, new_n137_})
2'b01 : new_n1577_ = 1'b1;
default : new_n1577_ = 1'b0;
endcase
casez ({new_n83_, new_n137_})
2'b01 : new_n1578_ = 1'b1;
default : new_n1578_ = 1'b0;
endcase
casez ({v[2], new_n141_})
2'b11 : new_n1579_ = 1'b1;
default : new_n1579_ = 1'b0;
endcase
casez ({y[1], new_n141_})
2'b11 : new_n1580_ = 1'b1;
default : new_n1580_ = 1'b0;
endcase
casez ({new_n81_, new_n141_})
2'b01 : new_n1581_ = 1'b1;
default : new_n1581_ = 1'b0;
endcase
casez ({new_n231_, new_n257_})
2'b11 : new_n1582_ = 1'b1;
default : new_n1582_ = 1'b0;
endcase
casez ({v[2], new_n147_})
2'b11 : new_n1583_ = 1'b1;
default : new_n1583_ = 1'b0;
endcase
casez ({new_n144_, new_n148_})
2'b11 : new_n1584_ = 1'b1;
default : new_n1584_ = 1'b0;
endcase
casez ({new_n118_, new_n151_})
2'b11 : new_n1585_ = 1'b1;
default : new_n1585_ = 1'b0;
endcase
casez ({new_n131_, new_n151_})
2'b11 : new_n1586_ = 1'b1;
default : new_n1586_ = 1'b0;
endcase
casez ({new_n151_, new_n153_})
2'b11 : new_n1587_ = 1'b1;
default : new_n1587_ = 1'b0;
endcase
casez ({new_n182_, new_n531_})
2'b11 : new_n1588_ = 1'b1;
default : new_n1588_ = 1'b0;
endcase
casez ({new_n104_, new_n275_})
2'b11 : new_n1589_ = 1'b1;
default : new_n1589_ = 1'b0;
endcase
casez ({new_n151_, new_n275_})
2'b11 : new_n1590_ = 1'b1;
default : new_n1590_ = 1'b0;
endcase
casez ({new_n148_, new_n160_})
2'b11 : new_n1591_ = 1'b1;
default : new_n1591_ = 1'b0;
endcase
casez ({new_n155_, new_n160_})
2'b11 : new_n1592_ = 1'b1;
default : new_n1592_ = 1'b0;
endcase
casez ({new_n155_, new_n162_})
2'b11 : new_n1593_ = 1'b1;
default : new_n1593_ = 1'b0;
endcase
casez ({new_n118_, new_n284_})
2'b11 : new_n1594_ = 1'b1;
default : new_n1594_ = 1'b0;
endcase
casez ({new_n115_, new_n166_})
2'b11 : new_n1595_ = 1'b1;
default : new_n1595_ = 1'b0;
endcase
casez ({new_n139_, new_n166_})
2'b11 : new_n1596_ = 1'b1;
default : new_n1596_ = 1'b0;
endcase
casez ({new_n154_, new_n166_})
2'b11 : new_n1597_ = 1'b1;
default : new_n1597_ = 1'b0;
endcase
casez ({new_n123_, new_n287_})
2'b11 : new_n1598_ = 1'b1;
default : new_n1598_ = 1'b0;
endcase
casez ({new_n166_, new_n169_})
2'b11 : new_n1599_ = 1'b1;
default : new_n1599_ = 1'b0;
endcase
casez ({new_n191_, new_n299_})
2'b11 : new_n1600_ = 1'b1;
default : new_n1600_ = 1'b0;
endcase
casez ({new_n162_, new_n174_})
2'b11 : new_n1601_ = 1'b1;
default : new_n1601_ = 1'b0;
endcase
casez ({new_n115_, new_n174_})
2'b11 : new_n1602_ = 1'b1;
default : new_n1602_ = 1'b0;
endcase
casez ({new_n142_, new_n174_})
2'b11 : new_n1603_ = 1'b1;
default : new_n1603_ = 1'b0;
endcase
casez ({new_n150_, new_n176_})
2'b11 : new_n1604_ = 1'b1;
default : new_n1604_ = 1'b0;
endcase
casez ({new_n94_, new_n180_})
2'b11 : new_n1605_ = 1'b1;
default : new_n1605_ = 1'b0;
endcase
casez ({new_n191_, new_n328_})
2'b11 : new_n1606_ = 1'b1;
default : new_n1606_ = 1'b0;
endcase
casez ({new_n115_, new_n187_})
2'b11 : new_n1607_ = 1'b1;
default : new_n1607_ = 1'b0;
endcase
casez ({new_n118_, new_n192_})
2'b11 : new_n1608_ = 1'b1;
default : new_n1608_ = 1'b0;
endcase
casez ({new_n139_, new_n192_})
2'b11 : new_n1609_ = 1'b1;
default : new_n1609_ = 1'b0;
endcase
casez ({u[1], new_n194_})
2'b11 : new_n1610_ = 1'b1;
default : new_n1610_ = 1'b0;
endcase
casez ({new_n94_, new_n194_})
2'b11 : new_n1611_ = 1'b1;
default : new_n1611_ = 1'b0;
endcase
casez ({new_n139_, new_n200_})
2'b11 : new_n1612_ = 1'b1;
default : new_n1612_ = 1'b0;
endcase
casez ({y[1], new_n357_})
2'b01 : new_n1613_ = 1'b1;
default : new_n1613_ = 1'b0;
endcase
casez ({new_n4616_, new_n95_, new_n940_})
3'b1?? : new_n1614_ = 1'b1;
3'b?11 : new_n1614_ = 1'b1;
default : new_n1614_ = 1'b0;
endcase
casez ({new_n131_, new_n208_})
2'b11 : new_n1615_ = 1'b1;
default : new_n1615_ = 1'b0;
endcase
casez ({new_n151_, new_n209_})
2'b11 : new_n1616_ = 1'b1;
default : new_n1616_ = 1'b0;
endcase
casez ({new_n182_, new_n211_})
2'b11 : new_n1617_ = 1'b1;
default : new_n1617_ = 1'b0;
endcase
casez ({new_n139_, new_n385_})
2'b11 : new_n1618_ = 1'b1;
default : new_n1618_ = 1'b0;
endcase
casez ({new_n93_, new_n204_})
2'b11 : new_n1619_ = 1'b1;
default : new_n1619_ = 1'b0;
endcase
casez ({v[1], new_n107_})
2'b10 : new_n1620_ = 1'b1;
default : new_n1620_ = 1'b0;
endcase
casez ({new_n167_, new_n219_})
2'b11 : new_n1621_ = 1'b1;
default : new_n1621_ = 1'b0;
endcase
casez ({new_n97_, new_n220_})
2'b11 : new_n1622_ = 1'b1;
default : new_n1622_ = 1'b0;
endcase
casez ({new_n94_, new_n219_})
2'b11 : new_n1623_ = 1'b1;
default : new_n1623_ = 1'b0;
endcase
casez ({new_n191_, new_n411_})
2'b11 : new_n1624_ = 1'b1;
default : new_n1624_ = 1'b0;
endcase
casez ({y[2], new_n222_})
2'b01 : new_n1625_ = 1'b1;
default : new_n1625_ = 1'b0;
endcase
casez ({new_n88_, new_n116_})
2'b01 : new_n1626_ = 1'b1;
default : new_n1626_ = 1'b0;
endcase
casez ({new_n118_, new_n230_})
2'b11 : new_n1627_ = 1'b1;
default : new_n1627_ = 1'b0;
endcase
casez ({new_n142_, new_n235_})
2'b11 : new_n1628_ = 1'b1;
default : new_n1628_ = 1'b0;
endcase
casez ({v[2], new_n128_})
2'b11 : new_n1629_ = 1'b1;
default : new_n1629_ = 1'b0;
endcase
casez ({new_n85_, new_n241_})
2'b11 : new_n1630_ = 1'b1;
default : new_n1630_ = 1'b0;
endcase
casez ({new_n103_, new_n243_})
2'b11 : new_n1631_ = 1'b1;
default : new_n1631_ = 1'b0;
endcase
casez ({new_n131_, new_n476_})
2'b11 : new_n1632_ = 1'b1;
default : new_n1632_ = 1'b0;
endcase
casez ({y[2], new_n145_})
2'b11 : new_n1633_ = 1'b1;
default : new_n1633_ = 1'b0;
endcase
casez ({v[1], new_n152_})
2'b01 : new_n1634_ = 1'b1;
default : new_n1634_ = 1'b0;
endcase
casez ({x[2], new_n154_})
2'b11 : new_n1635_ = 1'b1;
default : new_n1635_ = 1'b0;
endcase
casez ({new_n93_, new_n158_})
2'b11 : new_n1636_ = 1'b1;
default : new_n1636_ = 1'b0;
endcase
casez ({x[1], new_n160_})
2'b11 : new_n1637_ = 1'b1;
default : new_n1637_ = 1'b0;
endcase
casez ({new_n80_, new_n161_})
2'b11 : new_n1638_ = 1'b1;
default : new_n1638_ = 1'b0;
endcase
casez ({v[2], new_n154_})
2'b01 : new_n1639_ = 1'b1;
default : new_n1639_ = 1'b0;
endcase
casez ({x[1], new_n192_})
2'b11 : new_n1640_ = 1'b1;
default : new_n1640_ = 1'b0;
endcase
casez ({x[2], new_n194_})
2'b01 : new_n1641_ = 1'b1;
default : new_n1641_ = 1'b0;
endcase
casez ({x[1], new_n210_})
2'b11 : new_n1642_ = 1'b1;
default : new_n1642_ = 1'b0;
endcase
casez ({new_n84_, new_n109_})
2'b10 : new_n1643_ = 1'b1;
default : new_n1643_ = 1'b0;
endcase
casez ({new_n107_, new_n223_})
2'b01 : new_n1644_ = 1'b1;
default : new_n1644_ = 1'b0;
endcase
casez ({x[2], new_n115_})
2'b01 : new_n1645_ = 1'b1;
default : new_n1645_ = 1'b0;
endcase
casez ({new_n85_, new_n118_})
2'b11 : new_n1646_ = 1'b1;
default : new_n1646_ = 1'b0;
endcase
casez ({x[2], new_n118_})
2'b11 : new_n1647_ = 1'b1;
default : new_n1647_ = 1'b0;
endcase
casez ({new_n83_, new_n123_})
2'b11 : new_n1648_ = 1'b1;
default : new_n1648_ = 1'b0;
endcase
casez ({x[2], new_n131_})
2'b01 : new_n1649_ = 1'b1;
default : new_n1649_ = 1'b0;
endcase
casez ({u[0], new_n133_})
2'b11 : new_n1650_ = 1'b1;
default : new_n1650_ = 1'b0;
endcase
casez ({new_n98_, new_n135_})
2'b11 : new_n1651_ = 1'b1;
default : new_n1651_ = 1'b0;
endcase
casez ({new_n89_, new_n137_})
2'b11 : new_n1652_ = 1'b1;
default : new_n1652_ = 1'b0;
endcase
casez ({new_n142_, new_n155_, new_n1143_})
3'b11? : new_n1653_ = 1'b1;
3'b??1 : new_n1653_ = 1'b1;
default : new_n1653_ = 1'b0;
endcase
casez ({new_n3526_, new_n1146_})
2'b1? : new_n1654_ = 1'b1;
2'b?1 : new_n1654_ = 1'b1;
default : new_n1654_ = 1'b0;
endcase
casez ({new_n177_, new_n212_, new_n777_})
3'b11? : new_n1655_ = 1'b1;
3'b??1 : new_n1655_ = 1'b1;
default : new_n1655_ = 1'b0;
endcase
casez ({new_n189_, new_n305_, new_n1153_})
3'b11? : new_n1656_ = 1'b1;
3'b??1 : new_n1656_ = 1'b1;
default : new_n1656_ = 1'b0;
endcase
casez ({new_n4645_, new_n1155_})
2'b1? : new_n1657_ = 1'b1;
2'b?1 : new_n1657_ = 1'b1;
default : new_n1657_ = 1'b0;
endcase
casez ({new_n3495_, new_n1161_})
2'b1? : new_n1658_ = 1'b1;
2'b?1 : new_n1658_ = 1'b1;
default : new_n1658_ = 1'b0;
endcase
casez ({new_n194_, new_n764_, new_n784_})
3'b11? : new_n1659_ = 1'b1;
3'b??1 : new_n1659_ = 1'b1;
default : new_n1659_ = 1'b0;
endcase
casez ({new_n3326_, new_n1163_})
2'b1? : new_n1660_ = 1'b1;
2'b?1 : new_n1660_ = 1'b1;
default : new_n1660_ = 1'b0;
endcase
casez ({new_n3456_, new_n1167_})
2'b1? : new_n1661_ = 1'b1;
2'b?1 : new_n1661_ = 1'b1;
default : new_n1661_ = 1'b0;
endcase
casez ({new_n83_, new_n500_, new_n1176_})
3'b11? : new_n1662_ = 1'b1;
3'b??1 : new_n1662_ = 1'b1;
default : new_n1662_ = 1'b0;
endcase
casez ({new_n2579_, new_n543_})
2'b1? : new_n1663_ = 1'b1;
2'b?1 : new_n1663_ = 1'b1;
default : new_n1663_ = 1'b0;
endcase
casez ({new_n131_, new_n199_, new_n857_})
3'b11? : new_n1664_ = 1'b1;
3'b??1 : new_n1664_ = 1'b1;
default : new_n1664_ = 1'b0;
endcase
casez ({new_n4642_, new_n858_})
2'b1? : new_n1665_ = 1'b1;
2'b?1 : new_n1665_ = 1'b1;
default : new_n1665_ = 1'b0;
endcase
casez ({new_n150_, new_n254_, new_n295_})
3'b11? : new_n1666_ = 1'b1;
3'b??1 : new_n1666_ = 1'b1;
default : new_n1666_ = 1'b0;
endcase
casez ({new_n2502_, new_n871_})
2'b1? : new_n1667_ = 1'b1;
2'b?1 : new_n1667_ = 1'b1;
default : new_n1667_ = 1'b0;
endcase
casez ({new_n2726_, new_n871_})
2'b1? : new_n1668_ = 1'b1;
2'b?1 : new_n1668_ = 1'b1;
default : new_n1668_ = 1'b0;
endcase
casez ({new_n2137_, new_n1365_})
2'b1? : new_n1669_ = 1'b1;
2'b?1 : new_n1669_ = 1'b1;
default : new_n1669_ = 1'b0;
endcase
casez ({new_n2810_, new_n1380_})
2'b1? : new_n1670_ = 1'b1;
2'b?1 : new_n1670_ = 1'b1;
default : new_n1670_ = 1'b0;
endcase
casez ({new_n435_, new_n1390_})
2'b00 : new_n1671_ = 1'b1;
default : new_n1671_ = 1'b0;
endcase
casez ({new_n4646_, new_n384_})
2'b1? : new_n1672_ = 1'b1;
2'b?1 : new_n1672_ = 1'b1;
default : new_n1672_ = 1'b0;
endcase
casez ({new_n160_, new_n244_, new_n937_})
3'b11? : new_n1673_ = 1'b1;
3'b??1 : new_n1673_ = 1'b1;
default : new_n1673_ = 1'b0;
endcase
casez ({u[0], new_n340_, new_n620_})
3'b01? : new_n1674_ = 1'b1;
3'b??1 : new_n1674_ = 1'b1;
default : new_n1674_ = 1'b0;
endcase
casez ({new_n2680_, new_n938_})
2'b1? : new_n1675_ = 1'b1;
2'b?1 : new_n1675_ = 1'b1;
default : new_n1675_ = 1'b0;
endcase
casez ({u[0], new_n404_, new_n947_})
3'b01? : new_n1676_ = 1'b1;
3'b??1 : new_n1676_ = 1'b1;
default : new_n1676_ = 1'b0;
endcase
casez ({new_n2815_, new_n949_})
2'b1? : new_n1677_ = 1'b1;
2'b?1 : new_n1677_ = 1'b1;
default : new_n1677_ = 1'b0;
endcase
casez ({new_n86_, new_n207_, new_n952_})
3'b11? : new_n1678_ = 1'b1;
3'b??1 : new_n1678_ = 1'b1;
default : new_n1678_ = 1'b0;
endcase
casez ({new_n2712_, new_n956_})
2'b1? : new_n1679_ = 1'b1;
2'b?1 : new_n1679_ = 1'b1;
default : new_n1679_ = 1'b0;
endcase
casez ({new_n303_, new_n959_})
2'b00 : new_n1680_ = 1'b1;
default : new_n1680_ = 1'b0;
endcase
casez ({new_n2748_, new_n1010_})
2'b1? : new_n1681_ = 1'b1;
2'b?1 : new_n1681_ = 1'b1;
default : new_n1681_ = 1'b0;
endcase
casez ({new_n254_, new_n489_, new_n1017_})
3'b11? : new_n1682_ = 1'b1;
3'b??1 : new_n1682_ = 1'b1;
default : new_n1682_ = 1'b0;
endcase
casez ({new_n87_, new_n124_, new_n680_})
3'b11? : new_n1683_ = 1'b1;
3'b??1 : new_n1683_ = 1'b1;
default : new_n1683_ = 1'b0;
endcase
casez ({new_n85_, new_n1025_, new_n419_})
3'b01? : new_n1684_ = 1'b1;
3'b??1 : new_n1684_ = 1'b1;
default : new_n1684_ = 1'b0;
endcase
casez ({v[2], new_n483_, new_n1036_})
3'b11? : new_n1685_ = 1'b1;
3'b??1 : new_n1685_ = 1'b1;
default : new_n1685_ = 1'b0;
endcase
casez ({v[1], new_n478_, new_n1041_})
3'b11? : new_n1686_ = 1'b1;
3'b??1 : new_n1686_ = 1'b1;
default : new_n1686_ = 1'b0;
endcase
casez ({new_n84_, new_n729_, new_n384_})
3'b01? : new_n1687_ = 1'b1;
3'b??1 : new_n1687_ = 1'b1;
default : new_n1687_ = 1'b0;
endcase
casez ({new_n98_, new_n1094_, new_n863_})
3'b11? : new_n1688_ = 1'b1;
3'b??1 : new_n1688_ = 1'b1;
default : new_n1688_ = 1'b0;
endcase
casez ({new_n153_, new_n530_, new_n1106_})
3'b11? : new_n1689_ = 1'b1;
3'b??1 : new_n1689_ = 1'b1;
default : new_n1689_ = 1'b0;
endcase
casez ({new_n2674_, new_n1109_})
2'b1? : new_n1690_ = 1'b1;
2'b?1 : new_n1690_ = 1'b1;
default : new_n1690_ = 1'b0;
endcase
casez ({new_n2684_, new_n1111_})
2'b1? : new_n1691_ = 1'b1;
2'b?1 : new_n1691_ = 1'b1;
default : new_n1691_ = 1'b0;
endcase
casez ({new_n82_, new_n741_, new_n601_})
3'b01? : new_n1692_ = 1'b1;
3'b??1 : new_n1692_ = 1'b1;
default : new_n1692_ = 1'b0;
endcase
casez ({new_n88_, new_n275_, new_n1112_})
3'b11? : new_n1693_ = 1'b1;
3'b??1 : new_n1693_ = 1'b1;
default : new_n1693_ = 1'b0;
endcase
casez ({new_n3338_, new_n1115_})
2'b1? : new_n1694_ = 1'b1;
2'b?1 : new_n1694_ = 1'b1;
default : new_n1694_ = 1'b0;
endcase
casez ({new_n89_, new_n118_, new_n745_})
3'b11? : new_n1695_ = 1'b1;
3'b??1 : new_n1695_ = 1'b1;
default : new_n1695_ = 1'b0;
endcase
casez ({new_n3550_, new_n1121_})
2'b1? : new_n1696_ = 1'b1;
2'b?1 : new_n1696_ = 1'b1;
default : new_n1696_ = 1'b0;
endcase
casez ({new_n3520_, new_n1123_})
2'b1? : new_n1697_ = 1'b1;
2'b?1 : new_n1697_ = 1'b1;
default : new_n1697_ = 1'b0;
endcase
casez ({new_n2730_, new_n1124_})
2'b1? : new_n1698_ = 1'b1;
2'b?1 : new_n1698_ = 1'b1;
default : new_n1698_ = 1'b0;
endcase
casez ({x[1], new_n200_, new_n1125_})
3'b01? : new_n1699_ = 1'b1;
3'b??1 : new_n1699_ = 1'b1;
default : new_n1699_ = 1'b0;
endcase
casez ({new_n2836_, new_n1135_})
2'b1? : new_n1700_ = 1'b1;
2'b?1 : new_n1700_ = 1'b1;
default : new_n1700_ = 1'b0;
endcase
casez ({new_n3343_, new_n1136_})
2'b1? : new_n1701_ = 1'b1;
2'b?1 : new_n1701_ = 1'b1;
default : new_n1701_ = 1'b0;
endcase
casez ({new_n456_, new_n484_})
2'b00 : new_n1702_ = 1'b1;
default : new_n1702_ = 1'b0;
endcase
casez ({new_n605_, new_n776_})
2'b00 : new_n1703_ = 1'b1;
default : new_n1703_ = 1'b0;
endcase
casez ({new_n405_, new_n502_})
2'b00 : new_n1704_ = 1'b1;
default : new_n1704_ = 1'b0;
endcase
casez ({new_n3547_, new_n800_})
2'b1? : new_n1705_ = 1'b1;
2'b?1 : new_n1705_ = 1'b1;
default : new_n1705_ = 1'b0;
endcase
casez ({new_n389_, new_n524_})
2'b00 : new_n1706_ = 1'b1;
default : new_n1706_ = 1'b0;
endcase
casez ({new_n2768_, new_n295_})
2'b1? : new_n1707_ = 1'b1;
2'b?1 : new_n1707_ = 1'b1;
default : new_n1707_ = 1'b0;
endcase
casez ({new_n4654_, new_n289_})
2'b1? : new_n1708_ = 1'b1;
2'b?1 : new_n1708_ = 1'b1;
default : new_n1708_ = 1'b0;
endcase
casez ({new_n189_, new_n458_})
2'b00 : new_n1709_ = 1'b1;
default : new_n1709_ = 1'b0;
endcase
casez ({new_n361_, new_n457_})
2'b00 : new_n1710_ = 1'b1;
default : new_n1710_ = 1'b0;
endcase
casez ({new_n504_, new_n752_})
2'b00 : new_n1711_ = 1'b1;
default : new_n1711_ = 1'b0;
endcase
casez ({new_n122_, new_n251_})
2'b11 : new_n1712_ = 1'b1;
default : new_n1712_ = 1'b0;
endcase
casez ({new_n95_, new_n483_})
2'b11 : new_n1713_ = 1'b1;
default : new_n1713_ = 1'b0;
endcase
casez ({new_n157_, new_n254_})
2'b11 : new_n1714_ = 1'b1;
default : new_n1714_ = 1'b0;
endcase
casez ({new_n96_, new_n517_})
2'b11 : new_n1715_ = 1'b1;
default : new_n1715_ = 1'b0;
endcase
casez ({new_n94_, new_n483_})
2'b11 : new_n1716_ = 1'b1;
default : new_n1716_ = 1'b0;
endcase
casez ({u[1], new_n271_})
2'b11 : new_n1717_ = 1'b1;
default : new_n1717_ = 1'b0;
endcase
casez ({new_n79_, new_n272_})
2'b11 : new_n1718_ = 1'b1;
default : new_n1718_ = 1'b0;
endcase
casez ({new_n175_, new_n273_})
2'b11 : new_n1719_ = 1'b1;
default : new_n1719_ = 1'b0;
endcase
casez ({new_n156_, new_n558_})
2'b11 : new_n1720_ = 1'b1;
default : new_n1720_ = 1'b0;
endcase
casez ({new_n96_, new_n294_})
2'b11 : new_n1721_ = 1'b1;
default : new_n1721_ = 1'b0;
endcase
casez ({y[2], new_n324_})
2'b01 : new_n1722_ = 1'b1;
default : new_n1722_ = 1'b0;
endcase
casez ({v[2], new_n329_})
2'b11 : new_n1723_ = 1'b1;
default : new_n1723_ = 1'b0;
endcase
casez ({new_n171_, new_n198_})
2'b11 : new_n1724_ = 1'b1;
default : new_n1724_ = 1'b0;
endcase
casez ({new_n104_, new_n353_})
2'b11 : new_n1725_ = 1'b1;
default : new_n1725_ = 1'b0;
endcase
casez ({new_n86_, new_n353_})
2'b11 : new_n1726_ = 1'b1;
default : new_n1726_ = 1'b0;
endcase
casez ({x[0], new_n366_})
2'b11 : new_n1727_ = 1'b1;
default : new_n1727_ = 1'b0;
endcase
casez ({u[1], new_n371_})
2'b11 : new_n1728_ = 1'b1;
default : new_n1728_ = 1'b0;
endcase
casez ({new_n85_, new_n377_})
2'b11 : new_n1729_ = 1'b1;
default : new_n1729_ = 1'b0;
endcase
casez ({new_n104_, new_n377_})
2'b11 : new_n1730_ = 1'b1;
default : new_n1730_ = 1'b0;
endcase
casez ({new_n106_, new_n214_})
2'b11 : new_n1731_ = 1'b1;
default : new_n1731_ = 1'b0;
endcase
casez ({new_n86_, new_n389_})
2'b11 : new_n1732_ = 1'b1;
default : new_n1732_ = 1'b0;
endcase
casez ({new_n97_, new_n394_})
2'b10 : new_n1733_ = 1'b1;
default : new_n1733_ = 1'b0;
endcase
casez ({new_n223_, new_n398_})
2'b11 : new_n1734_ = 1'b1;
default : new_n1734_ = 1'b0;
endcase
casez ({new_n191_, new_n398_})
2'b11 : new_n1735_ = 1'b1;
default : new_n1735_ = 1'b0;
endcase
casez ({v[0], new_n397_})
2'b11 : new_n1736_ = 1'b1;
default : new_n1736_ = 1'b0;
endcase
casez ({x[0], new_n404_})
2'b11 : new_n1737_ = 1'b1;
default : new_n1737_ = 1'b0;
endcase
casez ({u[0], new_n407_})
2'b01 : new_n1738_ = 1'b1;
default : new_n1738_ = 1'b0;
endcase
casez ({y[0], new_n408_})
2'b11 : new_n1739_ = 1'b1;
default : new_n1739_ = 1'b0;
endcase
casez ({y[0], new_n421_})
2'b11 : new_n1740_ = 1'b1;
default : new_n1740_ = 1'b0;
endcase
casez ({new_n142_, new_n422_})
2'b11 : new_n1741_ = 1'b1;
default : new_n1741_ = 1'b0;
endcase
casez ({new_n148_, new_n420_})
2'b11 : new_n1742_ = 1'b1;
default : new_n1742_ = 1'b0;
endcase
casez ({u[0], new_n423_})
2'b11 : new_n1743_ = 1'b1;
default : new_n1743_ = 1'b0;
endcase
casez ({new_n114_, new_n124_})
2'b11 : new_n1744_ = 1'b1;
default : new_n1744_ = 1'b0;
endcase
casez ({new_n88_, new_n441_})
2'b11 : new_n1745_ = 1'b1;
default : new_n1745_ = 1'b0;
endcase
casez ({new_n122_, new_n237_})
2'b11 : new_n1746_ = 1'b1;
default : new_n1746_ = 1'b0;
endcase
casez ({new_n80_, new_n458_})
2'b11 : new_n1747_ = 1'b1;
default : new_n1747_ = 1'b0;
endcase
casez ({new_n79_, new_n280_})
2'b11 : new_n1748_ = 1'b1;
default : new_n1748_ = 1'b0;
endcase
casez ({new_n139_, new_n179_})
2'b11 : new_n1749_ = 1'b1;
default : new_n1749_ = 1'b0;
endcase
casez ({u[0], new_n181_})
2'b00 : new_n1750_ = 1'b1;
default : new_n1750_ = 1'b0;
endcase
casez ({new_n84_, new_n334_})
2'b11 : new_n1751_ = 1'b1;
default : new_n1751_ = 1'b0;
endcase
casez ({new_n97_, new_n360_})
2'b11 : new_n1752_ = 1'b1;
default : new_n1752_ = 1'b0;
endcase
casez ({new_n121_, new_n209_})
2'b11 : new_n1753_ = 1'b1;
default : new_n1753_ = 1'b0;
endcase
casez ({new_n101_, new_n390_})
2'b11 : new_n1754_ = 1'b1;
default : new_n1754_ = 1'b0;
endcase
casez ({new_n118_, new_n122_})
2'b11 : new_n1755_ = 1'b1;
default : new_n1755_ = 1'b0;
endcase
casez ({new_n2508_, new_n195_})
2'b1? : new_n1756_ = 1'b1;
2'b?1 : new_n1756_ = 1'b1;
default : new_n1756_ = 1'b0;
endcase
casez ({new_n83_, new_n333_, new_n296_})
3'b10? : new_n1757_ = 1'b1;
3'b??1 : new_n1757_ = 1'b1;
default : new_n1757_ = 1'b0;
endcase
casez ({new_n286_, new_n426_})
2'b00 : new_n1758_ = 1'b1;
default : new_n1758_ = 1'b0;
endcase
casez ({new_n2667_, new_n513_})
2'b1? : new_n1759_ = 1'b1;
2'b?1 : new_n1759_ = 1'b1;
default : new_n1759_ = 1'b0;
endcase
casez ({new_n3475_, new_n520_})
2'b1? : new_n1760_ = 1'b1;
2'b?1 : new_n1760_ = 1'b1;
default : new_n1760_ = 1'b0;
endcase
casez ({new_n3407_, new_n1202_})
2'b1? : new_n1761_ = 1'b1;
2'b?1 : new_n1761_ = 1'b1;
default : new_n1761_ = 1'b0;
endcase
casez ({new_n272_, new_n812_})
2'b00 : new_n1762_ = 1'b1;
default : new_n1762_ = 1'b0;
endcase
casez ({new_n153_, new_n246_, new_n814_})
3'b11? : new_n1763_ = 1'b1;
3'b??1 : new_n1763_ = 1'b1;
default : new_n1763_ = 1'b0;
endcase
casez ({new_n2598_, new_n1212_})
2'b1? : new_n1764_ = 1'b1;
2'b?1 : new_n1764_ = 1'b1;
default : new_n1764_ = 1'b0;
endcase
casez ({new_n188_, new_n539_})
2'b00 : new_n1765_ = 1'b1;
default : new_n1765_ = 1'b0;
endcase
casez ({new_n3555_, new_n839_})
2'b1? : new_n1766_ = 1'b1;
2'b?1 : new_n1766_ = 1'b1;
default : new_n1766_ = 1'b0;
endcase
casez ({y[2], new_n706_, new_n1304_})
3'b01? : new_n1767_ = 1'b1;
3'b??1 : new_n1767_ = 1'b1;
default : new_n1767_ = 1'b0;
endcase
casez ({new_n2653_, new_n568_})
2'b1? : new_n1768_ = 1'b1;
2'b?1 : new_n1768_ = 1'b1;
default : new_n1768_ = 1'b0;
endcase
casez ({new_n450_, new_n897_})
2'b00 : new_n1769_ = 1'b1;
default : new_n1769_ = 1'b0;
endcase
casez ({new_n3561_, new_n908_})
2'b1? : new_n1770_ = 1'b1;
2'b?1 : new_n1770_ = 1'b1;
default : new_n1770_ = 1'b0;
endcase
casez ({new_n168_, new_n444_, new_n658_})
3'b11? : new_n1771_ = 1'b1;
3'b??1 : new_n1771_ = 1'b1;
default : new_n1771_ = 1'b0;
endcase
casez ({new_n2636_, new_n662_})
2'b1? : new_n1772_ = 1'b1;
2'b?1 : new_n1772_ = 1'b1;
default : new_n1772_ = 1'b0;
endcase
casez ({y[2], new_n231_, new_n373_})
3'b01? : new_n1773_ = 1'b1;
3'b??1 : new_n1773_ = 1'b1;
default : new_n1773_ = 1'b0;
endcase
casez ({new_n3470_, new_n724_})
2'b1? : new_n1774_ = 1'b1;
2'b?1 : new_n1774_ = 1'b1;
default : new_n1774_ = 1'b0;
endcase
casez ({new_n197_, new_n739_})
2'b00 : new_n1775_ = 1'b1;
default : new_n1775_ = 1'b0;
endcase
casez ({new_n216_, new_n246_, new_n464_})
3'b11? : new_n1776_ = 1'b1;
3'b??1 : new_n1776_ = 1'b1;
default : new_n1776_ = 1'b0;
endcase
casez ({new_n3487_, new_n756_})
2'b1? : new_n1777_ = 1'b1;
2'b?1 : new_n1777_ = 1'b1;
default : new_n1777_ = 1'b0;
endcase
casez ({new_n2709_, new_n589_})
2'b1? : new_n1778_ = 1'b1;
2'b?1 : new_n1778_ = 1'b1;
default : new_n1778_ = 1'b0;
endcase
casez ({new_n103_, new_n888_, new_n1185_})
3'b11? : new_n1779_ = 1'b1;
3'b??1 : new_n1779_ = 1'b1;
default : new_n1779_ = 1'b0;
endcase
casez ({new_n2711_, new_n803_})
2'b1? : new_n1780_ = 1'b1;
2'b?1 : new_n1780_ = 1'b1;
default : new_n1780_ = 1'b0;
endcase
casez ({new_n214_, new_n813_, new_n1197_})
3'b11? : new_n1781_ = 1'b1;
3'b??1 : new_n1781_ = 1'b1;
default : new_n1781_ = 1'b0;
endcase
casez ({new_n2690_, new_n521_})
2'b1? : new_n1782_ = 1'b1;
2'b?1 : new_n1782_ = 1'b1;
default : new_n1782_ = 1'b0;
endcase
casez ({new_n168_, new_n531_, new_n547_})
3'b11? : new_n1783_ = 1'b1;
3'b??1 : new_n1783_ = 1'b1;
default : new_n1783_ = 1'b0;
endcase
casez ({new_n2824_, new_n882_})
2'b1? : new_n1784_ = 1'b1;
2'b?1 : new_n1784_ = 1'b1;
default : new_n1784_ = 1'b0;
endcase
casez ({new_n150_, new_n168_, new_n760_})
3'b11? : new_n1785_ = 1'b1;
3'b??1 : new_n1785_ = 1'b1;
default : new_n1785_ = 1'b0;
endcase
casez ({new_n117_, new_n257_})
2'b11 : new_n1786_ = 1'b1;
default : new_n1786_ = 1'b0;
endcase
casez ({new_n117_, new_n260_})
2'b11 : new_n1787_ = 1'b1;
default : new_n1787_ = 1'b0;
endcase
casez ({new_n149_, new_n563_})
2'b11 : new_n1788_ = 1'b1;
default : new_n1788_ = 1'b0;
endcase
casez ({new_n79_, new_n311_, new_n1077_})
3'b01? : new_n1789_ = 1'b1;
3'b??1 : new_n1789_ = 1'b1;
default : new_n1789_ = 1'b0;
endcase
casez ({new_n89_, new_n282_, new_n1086_})
3'b01? : new_n1790_ = 1'b1;
3'b??1 : new_n1790_ = 1'b1;
default : new_n1790_ = 1'b0;
endcase
casez ({new_n123_, new_n498_, new_n1244_})
3'b11? : new_n1791_ = 1'b1;
3'b??1 : new_n1791_ = 1'b1;
default : new_n1791_ = 1'b0;
endcase
casez ({new_n719_, new_n1062_, new_n1245_})
3'b11? : new_n1792_ = 1'b1;
3'b??1 : new_n1792_ = 1'b1;
default : new_n1792_ = 1'b0;
endcase
casez ({new_n281_, new_n617_, new_n918_})
3'b11? : new_n1793_ = 1'b1;
3'b??1 : new_n1793_ = 1'b1;
default : new_n1793_ = 1'b0;
endcase
casez ({new_n347_, new_n636_, new_n1252_})
3'b11? : new_n1794_ = 1'b1;
3'b??1 : new_n1794_ = 1'b1;
default : new_n1794_ = 1'b0;
endcase
casez ({new_n2821_, new_n920_})
2'b1? : new_n1795_ = 1'b1;
2'b?1 : new_n1795_ = 1'b1;
default : new_n1795_ = 1'b0;
endcase
casez ({u[2], v[1]})
2'b01 : new_n1796_ = 1'b1;
default : new_n1796_ = 1'b0;
endcase
casez ({u[1], new_n92_})
2'b11 : new_n1797_ = 1'b1;
default : new_n1797_ = 1'b0;
endcase
casez ({new_n88_, new_n95_})
2'b11 : new_n1798_ = 1'b1;
default : new_n1798_ = 1'b0;
endcase
casez ({new_n95_, new_n98_})
2'b11 : new_n1799_ = 1'b1;
default : new_n1799_ = 1'b0;
endcase
casez ({new_n95_, new_n101_})
2'b11 : new_n1800_ = 1'b1;
default : new_n1800_ = 1'b0;
endcase
casez ({v[0], new_n81_})
2'b10 : new_n1801_ = 1'b1;
default : new_n1801_ = 1'b0;
endcase
casez ({y[0], new_n81_})
2'b10 : new_n1802_ = 1'b1;
default : new_n1802_ = 1'b0;
endcase
casez ({new_n85_, new_n89_})
2'b01 : new_n1803_ = 1'b1;
default : new_n1803_ = 1'b0;
endcase
casez ({new_n79_, new_n98_})
2'b01 : new_n1804_ = 1'b1;
default : new_n1804_ = 1'b0;
endcase
casez ({new_n96_, new_n437_})
2'b11 : new_n1805_ = 1'b1;
default : new_n1805_ = 1'b0;
endcase
casez ({new_n98_, new_n234_})
2'b11 : new_n1806_ = 1'b1;
default : new_n1806_ = 1'b0;
endcase
casez ({new_n89_, new_n95_})
2'b11 : new_n1807_ = 1'b1;
default : new_n1807_ = 1'b0;
endcase
casez ({new_n81_, new_n98_})
2'b11 : new_n1808_ = 1'b1;
default : new_n1808_ = 1'b0;
endcase
casez ({new_n118_, new_n156_})
2'b00 : new_n1809_ = 1'b1;
default : new_n1809_ = 1'b0;
endcase
casez ({new_n174_, new_n300_})
2'b00 : new_n1810_ = 1'b1;
default : new_n1810_ = 1'b0;
endcase
casez ({new_n244_, new_n307_})
2'b00 : new_n1811_ = 1'b1;
default : new_n1811_ = 1'b0;
endcase
casez ({new_n299_, new_n313_})
2'b00 : new_n1812_ = 1'b1;
default : new_n1812_ = 1'b0;
endcase
casez ({new_n151_, new_n191_})
2'b00 : new_n1813_ = 1'b1;
default : new_n1813_ = 1'b0;
endcase
casez ({new_n177_, new_n192_})
2'b00 : new_n1814_ = 1'b1;
default : new_n1814_ = 1'b0;
endcase
casez ({new_n174_, new_n346_})
2'b00 : new_n1815_ = 1'b1;
default : new_n1815_ = 1'b0;
endcase
casez ({new_n176_, new_n204_})
2'b00 : new_n1816_ = 1'b1;
default : new_n1816_ = 1'b0;
endcase
casez ({new_n3416_, new_n234_, new_n565_})
3'b1?? : new_n1817_ = 1'b1;
3'b?11 : new_n1817_ = 1'b1;
default : new_n1817_ = 1'b0;
endcase
casez ({new_n160_, new_n210_})
2'b00 : new_n1818_ = 1'b1;
default : new_n1818_ = 1'b0;
endcase
casez ({new_n427_, new_n437_})
2'b00 : new_n1819_ = 1'b1;
default : new_n1819_ = 1'b0;
endcase
casez ({new_n293_, new_n1098_})
2'b00 : new_n1820_ = 1'b1;
default : new_n1820_ = 1'b0;
endcase
casez ({new_n127_, new_n240_})
2'b00 : new_n1821_ = 1'b1;
default : new_n1821_ = 1'b0;
endcase
casez ({new_n248_, new_n487_})
2'b11 : new_n1822_ = 1'b1;
default : new_n1822_ = 1'b0;
endcase
casez ({new_n223_, new_n489_})
2'b11 : new_n1823_ = 1'b1;
default : new_n1823_ = 1'b0;
endcase
casez ({new_n238_, new_n489_})
2'b11 : new_n1824_ = 1'b1;
default : new_n1824_ = 1'b0;
endcase
casez ({new_n137_, new_n257_})
2'b11 : new_n1825_ = 1'b1;
default : new_n1825_ = 1'b0;
endcase
casez ({new_n215_, new_n260_})
2'b11 : new_n1826_ = 1'b1;
default : new_n1826_ = 1'b0;
endcase
casez ({new_n204_, new_n262_})
2'b11 : new_n1827_ = 1'b1;
default : new_n1827_ = 1'b0;
endcase
casez ({new_n242_, new_n264_})
2'b11 : new_n1828_ = 1'b1;
default : new_n1828_ = 1'b0;
endcase
casez ({new_n210_, new_n508_})
2'b11 : new_n1829_ = 1'b1;
default : new_n1829_ = 1'b0;
endcase
casez ({new_n123_, new_n153_})
2'b11 : new_n1830_ = 1'b1;
default : new_n1830_ = 1'b0;
endcase
casez ({new_n251_, new_n273_})
2'b11 : new_n1831_ = 1'b1;
default : new_n1831_ = 1'b0;
endcase
casez ({new_n183_, new_n275_})
2'b11 : new_n1832_ = 1'b1;
default : new_n1832_ = 1'b0;
endcase
casez ({new_n150_, new_n281_})
2'b11 : new_n1833_ = 1'b1;
default : new_n1833_ = 1'b0;
endcase
casez ({new_n144_, new_n287_})
2'b11 : new_n1834_ = 1'b1;
default : new_n1834_ = 1'b0;
endcase
casez ({new_n82_, new_n169_})
2'b01 : new_n1835_ = 1'b1;
default : new_n1835_ = 1'b0;
endcase
casez ({new_n139_, new_n170_})
2'b11 : new_n1836_ = 1'b1;
default : new_n1836_ = 1'b0;
endcase
casez ({new_n241_, new_n301_})
2'b11 : new_n1837_ = 1'b1;
default : new_n1837_ = 1'b0;
endcase
casez ({new_n139_, new_n305_})
2'b11 : new_n1838_ = 1'b1;
default : new_n1838_ = 1'b0;
endcase
casez ({new_n187_, new_n309_})
2'b11 : new_n1839_ = 1'b1;
default : new_n1839_ = 1'b0;
endcase
casez ({new_n182_, new_n321_})
2'b11 : new_n1840_ = 1'b1;
default : new_n1840_ = 1'b0;
endcase
casez ({new_n144_, new_n328_})
2'b11 : new_n1841_ = 1'b1;
default : new_n1841_ = 1'b0;
endcase
casez ({new_n189_, new_n328_})
2'b11 : new_n1842_ = 1'b1;
default : new_n1842_ = 1'b0;
endcase
casez ({new_n78_, new_n924_})
2'b11 : new_n1843_ = 1'b1;
default : new_n1843_ = 1'b0;
endcase
casez ({new_n2849_, new_n4635_})
2'b1? : new_n1844_ = 1'b1;
2'b?1 : new_n1844_ = 1'b1;
default : new_n1844_ = 1'b0;
endcase
casez ({new_n169_, new_n190_})
2'b11 : new_n1845_ = 1'b1;
default : new_n1845_ = 1'b0;
endcase
casez ({new_n196_, new_n338_})
2'b11 : new_n1846_ = 1'b1;
default : new_n1846_ = 1'b0;
endcase
casez ({new_n139_, new_n196_})
2'b11 : new_n1847_ = 1'b1;
default : new_n1847_ = 1'b0;
endcase
casez ({u[1], new_n343_})
2'b11 : new_n1848_ = 1'b1;
default : new_n1848_ = 1'b0;
endcase
casez ({new_n222_, new_n344_})
2'b11 : new_n1849_ = 1'b1;
default : new_n1849_ = 1'b0;
endcase
casez ({new_n93_, new_n200_})
2'b01 : new_n1850_ = 1'b1;
default : new_n1850_ = 1'b0;
endcase
casez ({new_n90_, new_n654_})
2'b11 : new_n1851_ = 1'b1;
default : new_n1851_ = 1'b0;
endcase
casez ({new_n137_, new_n207_})
2'b11 : new_n1852_ = 1'b1;
default : new_n1852_ = 1'b0;
endcase
casez ({new_n144_, new_n207_})
2'b11 : new_n1853_ = 1'b1;
default : new_n1853_ = 1'b0;
endcase
casez ({new_n177_, new_n369_})
2'b11 : new_n1854_ = 1'b1;
default : new_n1854_ = 1'b0;
endcase
casez ({new_n196_, new_n369_})
2'b11 : new_n1855_ = 1'b1;
default : new_n1855_ = 1'b0;
endcase
casez ({new_n160_, new_n209_})
2'b11 : new_n1856_ = 1'b1;
default : new_n1856_ = 1'b0;
endcase
casez ({new_n170_, new_n209_})
2'b11 : new_n1857_ = 1'b1;
default : new_n1857_ = 1'b0;
endcase
casez ({new_n170_, new_n211_})
2'b11 : new_n1858_ = 1'b1;
default : new_n1858_ = 1'b0;
endcase
casez ({new_n196_, new_n216_})
2'b11 : new_n1859_ = 1'b1;
default : new_n1859_ = 1'b0;
endcase
casez ({new_n140_, new_n216_})
2'b11 : new_n1860_ = 1'b1;
default : new_n1860_ = 1'b0;
endcase
casez ({new_n204_, new_n220_})
2'b11 : new_n1861_ = 1'b1;
default : new_n1861_ = 1'b0;
endcase
casez ({new_n191_, new_n706_})
2'b11 : new_n1862_ = 1'b1;
default : new_n1862_ = 1'b0;
endcase
casez ({new_n131_, new_n223_})
2'b11 : new_n1863_ = 1'b1;
default : new_n1863_ = 1'b0;
endcase
casez ({new_n129_, new_n356_})
2'b11 : new_n1864_ = 1'b1;
default : new_n1864_ = 1'b0;
endcase
casez ({new_n166_, new_n432_})
2'b11 : new_n1865_ = 1'b1;
default : new_n1865_ = 1'b0;
endcase
casez ({new_n183_, new_n432_})
2'b11 : new_n1866_ = 1'b1;
default : new_n1866_ = 1'b0;
endcase
casez ({new_n81_, new_n130_})
2'b01 : new_n1867_ = 1'b1;
default : new_n1867_ = 1'b0;
endcase
casez ({new_n184_, new_n241_})
2'b11 : new_n1868_ = 1'b1;
default : new_n1868_ = 1'b0;
endcase
casez ({new_n176_, new_n243_})
2'b11 : new_n1869_ = 1'b1;
default : new_n1869_ = 1'b0;
endcase
casez ({new_n177_, new_n243_})
2'b11 : new_n1870_ = 1'b1;
default : new_n1870_ = 1'b0;
endcase
casez ({new_n81_, new_n136_})
2'b01 : new_n1871_ = 1'b1;
default : new_n1871_ = 1'b0;
endcase
casez ({new_n82_, new_n136_})
2'b01 : new_n1872_ = 1'b1;
default : new_n1872_ = 1'b0;
endcase
casez ({new_n191_, new_n247_})
2'b11 : new_n1873_ = 1'b1;
default : new_n1873_ = 1'b0;
endcase
casez ({new_n145_, new_n249_})
2'b11 : new_n1874_ = 1'b1;
default : new_n1874_ = 1'b0;
endcase
casez ({new_n167_, new_n249_})
2'b11 : new_n1875_ = 1'b1;
default : new_n1875_ = 1'b0;
endcase
casez ({new_n235_, new_n250_})
2'b11 : new_n1876_ = 1'b1;
default : new_n1876_ = 1'b0;
endcase
casez ({new_n170_, new_n250_})
2'b11 : new_n1877_ = 1'b1;
default : new_n1877_ = 1'b0;
endcase
casez ({new_n140_, new_n250_})
2'b11 : new_n1878_ = 1'b1;
default : new_n1878_ = 1'b0;
endcase
casez ({new_n153_, new_n251_})
2'b11 : new_n1879_ = 1'b1;
default : new_n1879_ = 1'b0;
endcase
casez ({v[1], new_n255_})
2'b11 : new_n1880_ = 1'b1;
default : new_n1880_ = 1'b0;
endcase
casez ({new_n96_, new_n262_})
2'b11 : new_n1881_ = 1'b1;
default : new_n1881_ = 1'b0;
endcase
casez ({y[1], new_n147_})
2'b11 : new_n1882_ = 1'b1;
default : new_n1882_ = 1'b0;
endcase
casez ({new_n81_, new_n150_})
2'b01 : new_n1883_ = 1'b1;
default : new_n1883_ = 1'b0;
endcase
casez ({new_n80_, new_n156_})
2'b01 : new_n1884_ = 1'b1;
default : new_n1884_ = 1'b0;
endcase
casez ({x[1], new_n158_})
2'b01 : new_n1885_ = 1'b1;
default : new_n1885_ = 1'b0;
endcase
casez ({new_n212_, new_n278_})
2'b11 : new_n1886_ = 1'b1;
default : new_n1886_ = 1'b0;
endcase
casez ({new_n115_, new_n284_})
2'b11 : new_n1887_ = 1'b1;
default : new_n1887_ = 1'b0;
endcase
casez ({new_n82_, new_n165_})
2'b01 : new_n1888_ = 1'b1;
default : new_n1888_ = 1'b0;
endcase
casez ({new_n77_, new_n165_})
2'b11 : new_n1889_ = 1'b1;
default : new_n1889_ = 1'b0;
endcase
casez ({new_n144_, new_n166_})
2'b11 : new_n1890_ = 1'b1;
default : new_n1890_ = 1'b0;
endcase
casez ({u[2], new_n167_})
2'b11 : new_n1891_ = 1'b1;
default : new_n1891_ = 1'b0;
endcase
casez ({new_n94_, new_n293_})
2'b11 : new_n1892_ = 1'b1;
default : new_n1892_ = 1'b0;
endcase
casez ({u[2], new_n170_})
2'b01 : new_n1893_ = 1'b1;
default : new_n1893_ = 1'b0;
endcase
casez ({new_n115_, new_n300_})
2'b11 : new_n1894_ = 1'b1;
default : new_n1894_ = 1'b0;
endcase
casez ({new_n148_, new_n174_})
2'b11 : new_n1895_ = 1'b1;
default : new_n1895_ = 1'b0;
endcase
casez ({new_n115_, new_n305_})
2'b11 : new_n1896_ = 1'b1;
default : new_n1896_ = 1'b0;
endcase
casez ({new_n153_, new_n306_})
2'b11 : new_n1897_ = 1'b1;
default : new_n1897_ = 1'b0;
endcase
casez ({new_n82_, new_n180_})
2'b11 : new_n1898_ = 1'b1;
default : new_n1898_ = 1'b0;
endcase
casez ({new_n123_, new_n317_})
2'b11 : new_n1899_ = 1'b1;
default : new_n1899_ = 1'b0;
endcase
casez ({new_n139_, new_n182_})
2'b11 : new_n1900_ = 1'b1;
default : new_n1900_ = 1'b0;
endcase
casez ({new_n115_, new_n184_})
2'b11 : new_n1901_ = 1'b1;
default : new_n1901_ = 1'b0;
endcase
casez ({new_n87_, new_n184_})
2'b01 : new_n1902_ = 1'b1;
default : new_n1902_ = 1'b0;
endcase
casez ({new_n208_, new_n328_})
2'b11 : new_n1903_ = 1'b1;
default : new_n1903_ = 1'b0;
endcase
casez ({new_n131_, new_n187_})
2'b11 : new_n1904_ = 1'b1;
default : new_n1904_ = 1'b0;
endcase
casez ({new_n248_, new_n332_})
2'b11 : new_n1905_ = 1'b1;
default : new_n1905_ = 1'b0;
endcase
casez ({new_n159_, new_n338_})
2'b11 : new_n1906_ = 1'b1;
default : new_n1906_ = 1'b0;
endcase
casez ({new_n140_, new_n192_})
2'b11 : new_n1907_ = 1'b1;
default : new_n1907_ = 1'b0;
endcase
casez ({new_n167_, new_n343_})
2'b11 : new_n1908_ = 1'b1;
default : new_n1908_ = 1'b0;
endcase
casez ({new_n80_, new_n200_})
2'b11 : new_n1909_ = 1'b1;
default : new_n1909_ = 1'b0;
endcase
casez ({new_n104_, new_n358_})
2'b11 : new_n1910_ = 1'b1;
default : new_n1910_ = 1'b0;
endcase
casez ({x[1], new_n204_})
2'b11 : new_n1911_ = 1'b1;
default : new_n1911_ = 1'b0;
endcase
casez ({new_n194_, new_n205_})
2'b11 : new_n1912_ = 1'b1;
default : new_n1912_ = 1'b0;
endcase
casez ({u[0], new_n206_})
2'b01 : new_n1913_ = 1'b1;
default : new_n1913_ = 1'b0;
endcase
casez ({new_n173_, new_n207_})
2'b11 : new_n1914_ = 1'b1;
default : new_n1914_ = 1'b0;
endcase
casez ({new_n159_, new_n207_})
2'b11 : new_n1915_ = 1'b1;
default : new_n1915_ = 1'b0;
endcase
casez ({new_n196_, new_n207_})
2'b11 : new_n1916_ = 1'b1;
default : new_n1916_ = 1'b0;
endcase
casez ({x[1], new_n208_})
2'b11 : new_n1917_ = 1'b1;
default : new_n1917_ = 1'b0;
endcase
casez ({new_n198_, new_n208_})
2'b11 : new_n1918_ = 1'b1;
default : new_n1918_ = 1'b0;
endcase
casez ({new_n145_, new_n207_})
2'b11 : new_n1919_ = 1'b1;
default : new_n1919_ = 1'b0;
endcase
casez ({new_n204_, new_n212_})
2'b11 : new_n1920_ = 1'b1;
default : new_n1920_ = 1'b0;
endcase
casez ({new_n158_, new_n212_})
2'b11 : new_n1921_ = 1'b1;
default : new_n1921_ = 1'b0;
endcase
casez ({new_n86_, new_n212_})
2'b11 : new_n1922_ = 1'b1;
default : new_n1922_ = 1'b0;
endcase
casez ({new_n190_, new_n214_})
2'b11 : new_n1923_ = 1'b1;
default : new_n1923_ = 1'b0;
endcase
casez ({new_n162_, new_n217_})
2'b11 : new_n1924_ = 1'b1;
default : new_n1924_ = 1'b0;
endcase
casez ({new_n83_, new_n218_})
2'b11 : new_n1925_ = 1'b1;
default : new_n1925_ = 1'b0;
endcase
casez ({new_n101_, new_n220_})
2'b11 : new_n1926_ = 1'b1;
default : new_n1926_ = 1'b0;
endcase
casez ({new_n148_, new_n221_})
2'b11 : new_n1927_ = 1'b1;
default : new_n1927_ = 1'b0;
endcase
casez ({new_n98_, new_n228_})
2'b11 : new_n1928_ = 1'b1;
default : new_n1928_ = 1'b0;
endcase
casez ({new_n154_, new_n230_})
2'b11 : new_n1929_ = 1'b1;
default : new_n1929_ = 1'b0;
endcase
casez ({new_n215_, new_n444_})
2'b11 : new_n1930_ = 1'b1;
default : new_n1930_ = 1'b0;
endcase
casez ({v[1], new_n129_})
2'b11 : new_n1931_ = 1'b1;
default : new_n1931_ = 1'b0;
endcase
casez ({v[1], new_n240_})
2'b11 : new_n1932_ = 1'b1;
default : new_n1932_ = 1'b0;
endcase
casez ({new_n118_, new_n242_})
2'b11 : new_n1933_ = 1'b1;
default : new_n1933_ = 1'b0;
endcase
casez ({new_n104_, new_n243_})
2'b11 : new_n1934_ = 1'b1;
default : new_n1934_ = 1'b0;
endcase
casez ({new_n109_, new_n133_})
2'b01 : new_n1935_ = 1'b1;
default : new_n1935_ = 1'b0;
endcase
casez ({new_n167_, new_n247_})
2'b11 : new_n1936_ = 1'b1;
default : new_n1936_ = 1'b0;
endcase
casez ({new_n103_, new_n140_})
2'b11 : new_n1937_ = 1'b1;
default : new_n1937_ = 1'b0;
endcase
casez ({new_n387_, new_n1173_, new_n4640_})
3'b11? : new_n1938_ = 1'b1;
3'b??1 : new_n1938_ = 1'b1;
default : new_n1938_ = 1'b0;
endcase
casez ({new_n86_, new_n142_})
2'b11 : new_n1939_ = 1'b1;
default : new_n1939_ = 1'b0;
endcase
casez ({y[2], new_n144_})
2'b11 : new_n1940_ = 1'b1;
default : new_n1940_ = 1'b0;
endcase
casez ({v[2], new_n147_})
2'b01 : new_n1941_ = 1'b1;
default : new_n1941_ = 1'b0;
endcase
casez ({u[1], new_n148_})
2'b01 : new_n1942_ = 1'b1;
default : new_n1942_ = 1'b0;
endcase
casez ({new_n85_, new_n154_})
2'b11 : new_n1943_ = 1'b1;
default : new_n1943_ = 1'b0;
endcase
casez ({y[2], new_n155_})
2'b11 : new_n1944_ = 1'b1;
default : new_n1944_ = 1'b0;
endcase
casez ({new_n83_, new_n155_})
2'b11 : new_n1945_ = 1'b1;
default : new_n1945_ = 1'b0;
endcase
casez ({new_n80_, new_n160_})
2'b11 : new_n1946_ = 1'b1;
default : new_n1946_ = 1'b0;
endcase
casez ({new_n97_, new_n163_})
2'b11 : new_n1947_ = 1'b1;
default : new_n1947_ = 1'b0;
endcase
casez ({v[1], new_n163_})
2'b01 : new_n1948_ = 1'b1;
default : new_n1948_ = 1'b0;
endcase
casez ({new_n93_, new_n182_})
2'b11 : new_n1949_ = 1'b1;
default : new_n1949_ = 1'b0;
endcase
casez ({new_n84_, new_n190_})
2'b11 : new_n1950_ = 1'b1;
default : new_n1950_ = 1'b0;
endcase
casez ({new_n80_, new_n192_})
2'b11 : new_n1951_ = 1'b1;
default : new_n1951_ = 1'b0;
endcase
casez ({x[2], new_n194_})
2'b11 : new_n1952_ = 1'b1;
default : new_n1952_ = 1'b0;
endcase
casez ({new_n127_, new_n183_})
2'b11 : new_n1953_ = 1'b1;
default : new_n1953_ = 1'b0;
endcase
casez ({new_n97_, new_n217_})
2'b11 : new_n1954_ = 1'b1;
default : new_n1954_ = 1'b0;
endcase
casez ({new_n84_, new_n107_})
2'b10 : new_n1955_ = 1'b1;
default : new_n1955_ = 1'b0;
endcase
casez ({y[2], new_n119_})
2'b01 : new_n1956_ = 1'b1;
default : new_n1956_ = 1'b0;
endcase
casez ({y[2], new_n119_})
2'b11 : new_n1957_ = 1'b1;
default : new_n1957_ = 1'b0;
endcase
casez ({u[2], new_n229_})
2'b11 : new_n1958_ = 1'b1;
default : new_n1958_ = 1'b0;
endcase
casez ({new_n101_, new_n127_})
2'b11 : new_n1959_ = 1'b1;
default : new_n1959_ = 1'b0;
endcase
casez ({new_n96_, new_n127_})
2'b11 : new_n1960_ = 1'b1;
default : new_n1960_ = 1'b0;
endcase
casez ({v[1], new_n135_})
2'b01 : new_n1961_ = 1'b1;
default : new_n1961_ = 1'b0;
endcase
casez ({u[2], new_n248_})
2'b11 : new_n1962_ = 1'b1;
default : new_n1962_ = 1'b0;
endcase
casez ({x[2], new_n139_})
2'b01 : new_n1963_ = 1'b1;
default : new_n1963_ = 1'b0;
endcase
casez ({u[1], new_n118_})
2'b01 : new_n1964_ = 1'b1;
default : new_n1964_ = 1'b0;
endcase
casez ({new_n155_, new_n171_})
2'b00 : new_n1965_ = 1'b1;
default : new_n1965_ = 1'b0;
endcase
casez ({new_n112_, new_n1144_, new_n4660_})
3'b11? : new_n1966_ = 1'b1;
3'b??1 : new_n1966_ = 1'b1;
default : new_n1966_ = 1'b0;
endcase
casez ({new_n196_, new_n780_, new_n422_, new_n1145_})
4'b11?? : new_n1967_ = 1'b1;
4'b??11 : new_n1967_ = 1'b1;
default : new_n1967_ = 1'b0;
endcase
casez ({new_n212_, new_n1907_, new_n228_, new_n384_})
4'b11?? : new_n1968_ = 1'b1;
4'b??11 : new_n1968_ = 1'b1;
default : new_n1968_ = 1'b0;
endcase
casez ({new_n577_, new_n1148_})
2'b00 : new_n1969_ = 1'b1;
default : new_n1969_ = 1'b0;
endcase
casez ({new_n81_, new_n785_, new_n175_, new_n1913_})
4'b11?? : new_n1970_ = 1'b1;
4'b??11 : new_n1970_ = 1'b1;
default : new_n1970_ = 1'b0;
endcase
casez ({new_n236_, new_n484_, new_n353_, new_n383_})
4'b11?? : new_n1971_ = 1'b1;
4'b??11 : new_n1971_ = 1'b1;
default : new_n1971_ = 1'b0;
endcase
casez ({new_n176_, new_n780_, new_n250_, new_n1150_})
4'b11?? : new_n1972_ = 1'b1;
4'b??11 : new_n1972_ = 1'b1;
default : new_n1972_ = 1'b0;
endcase
casez ({new_n4639_, new_n4581_})
2'b1? : new_n1973_ = 1'b1;
2'b?1 : new_n1973_ = 1'b1;
default : new_n1973_ = 1'b0;
endcase
casez ({new_n90_, new_n777_, new_n378_, new_n455_})
4'b11?? : new_n1974_ = 1'b1;
4'b??11 : new_n1974_ = 1'b1;
default : new_n1974_ = 1'b0;
endcase
casez ({new_n249_, new_n601_, new_n1029_, new_n1926_})
4'b11?? : new_n1975_ = 1'b1;
4'b??11 : new_n1975_ = 1'b1;
default : new_n1975_ = 1'b0;
endcase
casez ({new_n118_, new_n1153_, new_n120_, new_n680_})
4'b11?? : new_n1976_ = 1'b1;
4'b??11 : new_n1976_ = 1'b1;
default : new_n1976_ = 1'b0;
endcase
casez ({new_n208_, new_n778_, new_n278_, new_n617_})
4'b11?? : new_n1977_ = 1'b1;
4'b??11 : new_n1977_ = 1'b1;
default : new_n1977_ = 1'b0;
endcase
casez ({new_n144_, new_n740_, new_n4582_})
3'b11? : new_n1978_ = 1'b1;
3'b??1 : new_n1978_ = 1'b1;
default : new_n1978_ = 1'b0;
endcase
casez ({new_n154_, new_n1154_, new_n170_, new_n553_})
4'b11?? : new_n1979_ = 1'b1;
4'b??11 : new_n1979_ = 1'b1;
default : new_n1979_ = 1'b0;
endcase
casez ({new_n1108_, new_n1155_})
2'b00 : new_n1980_ = 1'b1;
default : new_n1980_ = 1'b0;
endcase
casez ({new_n286_, new_n484_, new_n330_, new_n1156_})
4'b11?? : new_n1981_ = 1'b1;
4'b??11 : new_n1981_ = 1'b1;
default : new_n1981_ = 1'b0;
endcase
casez ({new_n372_, new_n1156_, new_n441_, new_n632_})
4'b11?? : new_n1982_ = 1'b1;
4'b??11 : new_n1982_ = 1'b1;
default : new_n1982_ = 1'b0;
endcase
casez ({new_n311_, new_n1158_})
2'b00 : new_n1983_ = 1'b1;
default : new_n1983_ = 1'b0;
endcase
casez ({new_n145_, new_n1943_, new_n272_, new_n584_})
4'b11?? : new_n1984_ = 1'b1;
4'b??11 : new_n1984_ = 1'b1;
default : new_n1984_ = 1'b0;
endcase
casez ({new_n211_, new_n421_, new_n387_, new_n1160_})
4'b11?? : new_n1985_ = 1'b1;
4'b??11 : new_n1985_ = 1'b1;
default : new_n1985_ = 1'b0;
endcase
casez ({new_n240_, new_n677_, new_n336_, new_n1944_})
4'b11?? : new_n1986_ = 1'b1;
4'b??11 : new_n1986_ = 1'b1;
default : new_n1986_ = 1'b0;
endcase
casez ({new_n190_, new_n498_, new_n299_, new_n367_})
4'b11?? : new_n1987_ = 1'b1;
4'b??11 : new_n1987_ = 1'b1;
default : new_n1987_ = 1'b0;
endcase
casez ({new_n247_, new_n471_, new_n748_, new_n1957_})
4'b11?? : new_n1988_ = 1'b1;
4'b??11 : new_n1988_ = 1'b1;
default : new_n1988_ = 1'b0;
endcase
casez ({new_n95_, new_n785_, new_n310_, new_n505_})
4'b11?? : new_n1989_ = 1'b1;
4'b??11 : new_n1989_ = 1'b1;
default : new_n1989_ = 1'b0;
endcase
casez ({new_n202_, new_n964_, new_n280_, new_n1167_})
4'b11?? : new_n1990_ = 1'b1;
4'b??11 : new_n1990_ = 1'b1;
default : new_n1990_ = 1'b0;
endcase
casez ({new_n185_, new_n502_, new_n339_, new_n340_})
4'b11?? : new_n1991_ = 1'b1;
4'b??11 : new_n1991_ = 1'b1;
default : new_n1991_ = 1'b0;
endcase
casez ({new_n155_, new_n788_, new_n310_, new_n372_})
4'b11?? : new_n1992_ = 1'b1;
4'b??11 : new_n1992_ = 1'b1;
default : new_n1992_ = 1'b0;
endcase
casez ({new_n86_, new_n738_, new_n447_, new_n1172_})
4'b11?? : new_n1993_ = 1'b1;
4'b??11 : new_n1993_ = 1'b1;
default : new_n1993_ = 1'b0;
endcase
casez ({new_n132_, new_n367_, new_n215_, new_n789_})
4'b11?? : new_n1994_ = 1'b1;
4'b??11 : new_n1994_ = 1'b1;
default : new_n1994_ = 1'b0;
endcase
casez ({new_n247_, new_n944_, new_n4586_})
3'b11? : new_n1995_ = 1'b1;
3'b??1 : new_n1995_ = 1'b1;
default : new_n1995_ = 1'b0;
endcase
casez ({new_n166_, new_n1004_, new_n632_, new_n1175_})
4'b11?? : new_n1996_ = 1'b1;
4'b??11 : new_n1996_ = 1'b1;
default : new_n1996_ = 1'b0;
endcase
casez ({new_n1039_, new_n1177_})
2'b00 : new_n1997_ = 1'b1;
default : new_n1997_ = 1'b0;
endcase
casez ({new_n501_, new_n525_})
2'b00 : new_n1998_ = 1'b1;
default : new_n1998_ = 1'b0;
endcase
casez ({new_n323_, new_n525_})
2'b00 : new_n1999_ = 1'b1;
default : new_n1999_ = 1'b0;
endcase
casez ({new_n324_, new_n538_})
2'b00 : new_n2000_ = 1'b1;
default : new_n2000_ = 1'b0;
endcase
casez ({new_n404_, new_n540_})
2'b00 : new_n2001_ = 1'b1;
default : new_n2001_ = 1'b0;
endcase
casez ({new_n88_, new_n854_, new_n4665_})
3'b11? : new_n2002_ = 1'b1;
3'b??1 : new_n2002_ = 1'b1;
default : new_n2002_ = 1'b0;
endcase
casez ({new_n230_, new_n854_, new_n401_, new_n580_})
4'b11?? : new_n2003_ = 1'b1;
4'b??11 : new_n2003_ = 1'b1;
default : new_n2003_ = 1'b0;
endcase
casez ({new_n735_, new_n856_})
2'b00 : new_n2004_ = 1'b1;
default : new_n2004_ = 1'b0;
endcase
casez ({new_n94_, new_n859_, new_n121_, new_n367_})
4'b11?? : new_n2005_ = 1'b1;
4'b??11 : new_n2005_ = 1'b1;
default : new_n2005_ = 1'b0;
endcase
casez ({new_n237_, new_n860_, new_n267_, new_n384_})
4'b11?? : new_n2006_ = 1'b1;
4'b??11 : new_n2006_ = 1'b1;
default : new_n2006_ = 1'b0;
endcase
casez ({new_n157_, new_n382_, new_n267_, new_n862_})
4'b11?? : new_n2007_ = 1'b1;
4'b??11 : new_n2007_ = 1'b1;
default : new_n2007_ = 1'b0;
endcase
casez ({new_n142_, new_n631_, new_n330_, new_n863_})
4'b11?? : new_n2008_ = 1'b1;
4'b??11 : new_n2008_ = 1'b1;
default : new_n2008_ = 1'b0;
endcase
casez ({new_n127_, new_n367_, new_n372_, new_n863_})
4'b11?? : new_n2009_ = 1'b1;
4'b??11 : new_n2009_ = 1'b1;
default : new_n2009_ = 1'b0;
endcase
casez ({new_n175_, new_n423_, new_n219_, new_n865_})
4'b11?? : new_n2010_ = 1'b1;
4'b??11 : new_n2010_ = 1'b1;
default : new_n2010_ = 1'b0;
endcase
casez ({new_n98_, new_n867_, new_n160_, new_n311_})
4'b11?? : new_n2011_ = 1'b1;
4'b??11 : new_n2011_ = 1'b1;
default : new_n2011_ = 1'b0;
endcase
casez ({new_n265_, new_n872_})
2'b00 : new_n2012_ = 1'b1;
default : new_n2012_ = 1'b0;
endcase
casez ({new_n173_, new_n185_, new_n199_, new_n577_})
4'b11?? : new_n2013_ = 1'b1;
4'b??11 : new_n2013_ = 1'b1;
default : new_n2013_ = 1'b0;
endcase
casez ({new_n501_, new_n872_})
2'b00 : new_n2014_ = 1'b1;
default : new_n2014_ = 1'b0;
endcase
casez ({new_n169_, new_n1337_, new_n290_, new_n874_})
4'b11?? : new_n2015_ = 1'b1;
4'b??11 : new_n2015_ = 1'b1;
default : new_n2015_ = 1'b0;
endcase
casez ({new_n80_, new_n746_, new_n243_, new_n1337_})
4'b11?? : new_n2016_ = 1'b1;
4'b??11 : new_n2016_ = 1'b1;
default : new_n2016_ = 1'b0;
endcase
casez ({new_n747_, new_n873_})
2'b00 : new_n2017_ = 1'b1;
default : new_n2017_ = 1'b0;
endcase
casez ({new_n116_, new_n259_, new_n167_, new_n580_})
4'b11?? : new_n2018_ = 1'b1;
4'b??11 : new_n2018_ = 1'b1;
default : new_n2018_ = 1'b0;
endcase
casez ({new_n132_, new_n1346_, new_n241_, new_n678_})
4'b11?? : new_n2019_ = 1'b1;
4'b??11 : new_n2019_ = 1'b1;
default : new_n2019_ = 1'b0;
endcase
casez ({new_n157_, new_n858_, new_n225_, new_n1347_})
4'b11?? : new_n2020_ = 1'b1;
4'b??11 : new_n2020_ = 1'b1;
default : new_n2020_ = 1'b0;
endcase
casez ({new_n2844_, new_n4595_})
2'b1? : new_n2021_ = 1'b1;
2'b?1 : new_n2021_ = 1'b1;
default : new_n2021_ = 1'b0;
endcase
casez ({new_n638_, new_n1351_})
2'b00 : new_n2022_ = 1'b1;
default : new_n2022_ = 1'b0;
endcase
casez ({new_n176_, new_n861_, new_n205_, new_n1352_})
4'b11?? : new_n2023_ = 1'b1;
4'b??11 : new_n2023_ = 1'b1;
default : new_n2023_ = 1'b0;
endcase
casez ({new_n1040_, new_n1366_})
2'b00 : new_n2024_ = 1'b1;
default : new_n2024_ = 1'b0;
endcase
casez ({new_n228_, new_n779_, new_n447_, new_n1367_})
4'b11?? : new_n2025_ = 1'b1;
4'b??11 : new_n2025_ = 1'b1;
default : new_n2025_ = 1'b0;
endcase
casez ({new_n430_, new_n601_, new_n460_, new_n1367_})
4'b11?? : new_n2026_ = 1'b1;
4'b??11 : new_n2026_ = 1'b1;
default : new_n2026_ = 1'b0;
endcase
casez ({new_n190_, new_n556_, new_n384_, new_n597_})
4'b11?? : new_n2027_ = 1'b1;
4'b??11 : new_n2027_ = 1'b1;
default : new_n2027_ = 1'b0;
endcase
casez ({new_n1139_, new_n1368_})
2'b00 : new_n2028_ = 1'b1;
default : new_n2028_ = 1'b0;
endcase
casez ({new_n127_, new_n419_, new_n284_, new_n600_})
4'b11?? : new_n2029_ = 1'b1;
4'b??11 : new_n2029_ = 1'b1;
default : new_n2029_ = 1'b0;
endcase
casez ({new_n137_, new_n419_, new_n210_, new_n600_})
4'b11?? : new_n2030_ = 1'b1;
4'b??11 : new_n2030_ = 1'b1;
default : new_n2030_ = 1'b0;
endcase
casez ({new_n4628_, new_n301_, new_n1381_})
3'b1?? : new_n2031_ = 1'b1;
3'b?11 : new_n2031_ = 1'b1;
default : new_n2031_ = 1'b0;
endcase
casez ({new_n158_, new_n1391_, new_n171_, new_n1141_})
4'b11?? : new_n2032_ = 1'b1;
4'b??11 : new_n2032_ = 1'b1;
default : new_n2032_ = 1'b0;
endcase
casez ({new_n259_, new_n324_, new_n290_, new_n1392_})
4'b11?? : new_n2033_ = 1'b1;
4'b??11 : new_n2033_ = 1'b1;
default : new_n2033_ = 1'b0;
endcase
casez ({new_n378_, new_n965_, new_n504_, new_n1394_})
4'b11?? : new_n2034_ = 1'b1;
4'b??11 : new_n2034_ = 1'b1;
default : new_n2034_ = 1'b0;
endcase
casez ({new_n240_, new_n1014_, new_n336_, new_n1400_})
4'b11?? : new_n2035_ = 1'b1;
4'b??11 : new_n2035_ = 1'b1;
default : new_n2035_ = 1'b0;
endcase
casez ({new_n190_, new_n1401_, new_n252_, new_n1003_})
4'b11?? : new_n2036_ = 1'b1;
4'b??01 : new_n2036_ = 1'b1;
default : new_n2036_ = 1'b0;
endcase
casez ({new_n350_, new_n959_, new_n454_, new_n1403_})
4'b11?? : new_n2037_ = 1'b1;
4'b??11 : new_n2037_ = 1'b1;
default : new_n2037_ = 1'b0;
endcase
casez ({new_n124_, new_n750_, new_n199_, new_n938_})
4'b11?? : new_n2038_ = 1'b1;
4'b??11 : new_n2038_ = 1'b1;
default : new_n2038_ = 1'b0;
endcase
casez ({new_n423_, new_n939_})
2'b00 : new_n2039_ = 1'b1;
default : new_n2039_ = 1'b0;
endcase
casez ({new_n345_, new_n634_, new_n366_, new_n447_})
4'b11?? : new_n2040_ = 1'b1;
4'b??11 : new_n2040_ = 1'b1;
default : new_n2040_ = 1'b0;
endcase
casez ({new_n430_, new_n951_, new_n482_, new_n774_})
4'b11?? : new_n2041_ = 1'b1;
4'b??10 : new_n2041_ = 1'b1;
default : new_n2041_ = 1'b0;
endcase
casez ({new_n458_, new_n503_, new_n863_, new_n953_})
4'b11?? : new_n2042_ = 1'b1;
4'b??11 : new_n2042_ = 1'b1;
default : new_n2042_ = 1'b0;
endcase
casez ({new_n183_, new_n668_, new_n221_, new_n954_})
4'b11?? : new_n2043_ = 1'b1;
4'b??11 : new_n2043_ = 1'b1;
default : new_n2043_ = 1'b0;
endcase
casez ({new_n351_, new_n954_, new_n367_, new_n707_})
4'b11?? : new_n2044_ = 1'b1;
4'b??10 : new_n2044_ = 1'b1;
default : new_n2044_ = 1'b0;
endcase
casez ({new_n175_, new_n638_, new_n377_, new_n957_})
4'b11?? : new_n2045_ = 1'b1;
4'b??11 : new_n2045_ = 1'b1;
default : new_n2045_ = 1'b0;
endcase
casez ({new_n292_, new_n959_, new_n303_, new_n729_})
4'b11?? : new_n2046_ = 1'b1;
4'b??11 : new_n2046_ = 1'b1;
default : new_n2046_ = 1'b0;
endcase
casez ({new_n715_, new_n962_})
2'b00 : new_n2047_ = 1'b1;
default : new_n2047_ = 1'b0;
endcase
casez ({new_n955_, new_n962_})
2'b00 : new_n2048_ = 1'b1;
default : new_n2048_ = 1'b0;
endcase
casez ({new_n236_, new_n1546_})
2'b00 : new_n2049_ = 1'b1;
default : new_n2049_ = 1'b0;
endcase
casez ({new_n766_, new_n1556_, new_n1095_, new_n1355_})
4'b11?? : new_n2050_ = 1'b1;
4'b??11 : new_n2050_ = 1'b1;
default : new_n2050_ = 1'b0;
endcase
casez ({new_n1114_, new_n1558_})
2'b00 : new_n2051_ = 1'b1;
default : new_n2051_ = 1'b0;
endcase
casez ({new_n144_, new_n1043_, new_n191_, new_n1561_})
4'b11?? : new_n2052_ = 1'b1;
4'b??11 : new_n2052_ = 1'b1;
default : new_n2052_ = 1'b0;
endcase
casez ({new_n122_, new_n384_, new_n201_, new_n1562_})
4'b11?? : new_n2053_ = 1'b1;
4'b??11 : new_n2053_ = 1'b1;
default : new_n2053_ = 1'b0;
endcase
casez ({new_n218_, new_n1564_, new_n306_, new_n1116_})
4'b11?? : new_n2054_ = 1'b1;
4'b??11 : new_n2054_ = 1'b1;
default : new_n2054_ = 1'b0;
endcase
casez ({new_n1028_, new_n1565_})
2'b00 : new_n2055_ = 1'b1;
default : new_n2055_ = 1'b0;
endcase
casez ({new_n481_, new_n620_, new_n965_, new_n1579_})
4'b11?? : new_n2056_ = 1'b1;
4'b??11 : new_n2056_ = 1'b1;
default : new_n2056_ = 1'b0;
endcase
casez ({new_n255_, new_n1008_, new_n419_, new_n706_})
4'b11?? : new_n2057_ = 1'b1;
4'b??11 : new_n2057_ = 1'b1;
default : new_n2057_ = 1'b0;
endcase
casez ({new_n295_, new_n1009_})
2'b00 : new_n2058_ = 1'b1;
default : new_n2058_ = 1'b0;
endcase
casez ({new_n540_, new_n1009_})
2'b00 : new_n2059_ = 1'b1;
default : new_n2059_ = 1'b0;
endcase
casez ({new_n161_, new_n1011_, new_n176_, new_n668_})
4'b11?? : new_n2060_ = 1'b1;
4'b??11 : new_n2060_ = 1'b1;
default : new_n2060_ = 1'b0;
endcase
casez ({new_n963_, new_n1587_})
2'b00 : new_n2061_ = 1'b1;
default : new_n2061_ = 1'b0;
endcase
casez ({new_n946_, new_n1014_})
2'b00 : new_n2062_ = 1'b1;
default : new_n2062_ = 1'b0;
endcase
casez ({new_n167_, new_n1122_, new_n262_, new_n1591_})
4'b11?? : new_n2063_ = 1'b1;
4'b??11 : new_n2063_ = 1'b1;
default : new_n2063_ = 1'b0;
endcase
casez ({new_n1116_, new_n1594_})
2'b00 : new_n2064_ = 1'b1;
default : new_n2064_ = 1'b0;
endcase
casez ({new_n103_, new_n580_, new_n115_, new_n681_})
4'b11?? : new_n2065_ = 1'b1;
4'b??11 : new_n2065_ = 1'b1;
default : new_n2065_ = 1'b0;
endcase
casez ({new_n482_, new_n1018_})
2'b00 : new_n2066_ = 1'b1;
default : new_n2066_ = 1'b0;
endcase
casez ({new_n182_, new_n1020_})
2'b00 : new_n2067_ = 1'b1;
default : new_n2067_ = 1'b0;
endcase
casez ({new_n1020_, new_n1023_})
2'b00 : new_n2068_ = 1'b1;
default : new_n2068_ = 1'b0;
endcase
casez ({new_n956_, new_n1023_})
2'b00 : new_n2069_ = 1'b1;
default : new_n2069_ = 1'b0;
endcase
casez ({new_n4623_, new_n299_, new_n1618_})
3'b1?? : new_n2070_ = 1'b1;
3'b?11 : new_n2070_ = 1'b1;
default : new_n2070_ = 1'b0;
endcase
casez ({new_n202_, new_n956_, new_n239_, new_n1621_})
4'b11?? : new_n2071_ = 1'b1;
4'b??11 : new_n2071_ = 1'b1;
default : new_n2071_ = 1'b0;
endcase
casez ({new_n745_, new_n1627_})
2'b00 : new_n2072_ = 1'b1;
default : new_n2072_ = 1'b0;
endcase
casez ({new_n267_, new_n367_, new_n391_, new_n1644_})
4'b11?? : new_n2073_ = 1'b1;
4'b??11 : new_n2073_ = 1'b1;
default : new_n2073_ = 1'b0;
endcase
casez ({new_n248_, new_n938_, new_n372_, new_n1647_})
4'b11?? : new_n2074_ = 1'b1;
4'b??11 : new_n2074_ = 1'b1;
default : new_n2074_ = 1'b0;
endcase
casez ({new_n737_, new_n1043_})
2'b00 : new_n2075_ = 1'b1;
default : new_n2075_ = 1'b0;
endcase
casez ({new_n638_, new_n1046_})
2'b00 : new_n2076_ = 1'b1;
default : new_n2076_ = 1'b0;
endcase
casez ({new_n207_, new_n951_, new_n447_, new_n1047_})
4'b11?? : new_n2077_ = 1'b1;
4'b??11 : new_n2077_ = 1'b1;
default : new_n2077_ = 1'b0;
endcase
casez ({new_n311_, new_n714_, new_n497_, new_n683_})
4'b11?? : new_n2078_ = 1'b1;
4'b??11 : new_n2078_ = 1'b1;
default : new_n2078_ = 1'b0;
endcase
casez ({new_n126_, new_n716_})
2'b00 : new_n2079_ = 1'b1;
default : new_n2079_ = 1'b0;
endcase
casez ({new_n290_, new_n423_, new_n313_, new_n367_})
4'b11?? : new_n2080_ = 1'b1;
4'b??11 : new_n2080_ = 1'b1;
default : new_n2080_ = 1'b0;
endcase
casez ({new_n454_, new_n734_})
2'b00 : new_n2081_ = 1'b1;
default : new_n2081_ = 1'b0;
endcase
casez ({new_n244_, new_n994_, new_n866_, new_n1095_})
4'b11?? : new_n2082_ = 1'b1;
4'b??11 : new_n2082_ = 1'b1;
default : new_n2082_ = 1'b0;
endcase
casez ({new_n339_, new_n749_, new_n958_, new_n1099_})
4'b11?? : new_n2083_ = 1'b1;
4'b??11 : new_n2083_ = 1'b1;
default : new_n2083_ = 1'b0;
endcase
casez ({new_n342_, new_n384_, new_n501_, new_n1102_})
4'b11?? : new_n2084_ = 1'b1;
4'b??11 : new_n2084_ = 1'b1;
default : new_n2084_ = 1'b0;
endcase
casez ({new_n200_, new_n577_, new_n267_, new_n737_})
4'b11?? : new_n2085_ = 1'b1;
4'b??11 : new_n2085_ = 1'b1;
default : new_n2085_ = 1'b0;
endcase
casez ({new_n179_, new_n798_, new_n634_, new_n1107_})
4'b11?? : new_n2086_ = 1'b1;
4'b??11 : new_n2086_ = 1'b1;
default : new_n2086_ = 1'b0;
endcase
casez ({new_n131_, new_n1827_, new_n293_, new_n1044_})
4'b11?? : new_n2087_ = 1'b1;
4'b??11 : new_n2087_ = 1'b1;
default : new_n2087_ = 1'b0;
endcase
casez ({new_n196_, new_n1834_, new_n211_, new_n937_})
4'b11?? : new_n2088_ = 1'b1;
4'b??11 : new_n2088_ = 1'b1;
default : new_n2088_ = 1'b0;
endcase
casez ({new_n329_, new_n1835_, new_n579_, new_n768_})
4'b11?? : new_n2089_ = 1'b1;
4'b??11 : new_n2089_ = 1'b1;
default : new_n2089_ = 1'b0;
endcase
casez ({new_n552_, new_n747_})
2'b00 : new_n2090_ = 1'b1;
default : new_n2090_ = 1'b0;
endcase
casez ({new_n265_, new_n747_})
2'b00 : new_n2091_ = 1'b1;
default : new_n2091_ = 1'b0;
endcase
casez ({new_n113_, new_n540_, new_n305_, new_n1127_})
4'b11?? : new_n2092_ = 1'b1;
4'b??11 : new_n2092_ = 1'b1;
default : new_n2092_ = 1'b0;
endcase
casez ({new_n151_, new_n1864_, new_n264_, new_n1592_})
4'b11?? : new_n2093_ = 1'b1;
4'b??11 : new_n2093_ = 1'b1;
default : new_n2093_ = 1'b0;
endcase
casez ({new_n1015_, new_n1130_})
2'b00 : new_n2094_ = 1'b1;
default : new_n2094_ = 1'b0;
endcase
casez ({new_n857_, new_n1130_})
2'b00 : new_n2095_ = 1'b1;
default : new_n2095_ = 1'b0;
endcase
casez ({new_n218_, new_n1868_, new_n504_, new_n683_})
4'b11?? : new_n2096_ = 1'b1;
4'b??11 : new_n2096_ = 1'b1;
default : new_n2096_ = 1'b0;
endcase
casez ({u[1], new_n1878_, new_n103_, new_n1358_})
4'b01?? : new_n2097_ = 1'b1;
4'b??11 : new_n2097_ = 1'b1;
default : new_n2097_ = 1'b0;
endcase
casez ({new_n395_, new_n1883_, new_n450_, new_n1016_})
4'b11?? : new_n2098_ = 1'b1;
4'b??11 : new_n2098_ = 1'b1;
default : new_n2098_ = 1'b0;
endcase
casez ({new_n330_, new_n868_, new_n345_, new_n1888_})
4'b11?? : new_n2099_ = 1'b1;
4'b??11 : new_n2099_ = 1'b1;
default : new_n2099_ = 1'b0;
endcase
casez ({new_n225_, new_n1021_, new_n1402_, new_n1889_})
4'b11?? : new_n2100_ = 1'b1;
4'b??11 : new_n2100_ = 1'b1;
default : new_n2100_ = 1'b0;
endcase
casez ({new_n862_, new_n1141_})
2'b00 : new_n2101_ = 1'b1;
default : new_n2101_ = 1'b0;
endcase
casez ({new_n157_, new_n495_})
2'b00 : new_n2102_ = 1'b1;
default : new_n2102_ = 1'b0;
endcase
casez ({new_n238_, new_n795_})
2'b00 : new_n2103_ = 1'b1;
default : new_n2103_ = 1'b0;
endcase
casez ({new_n424_, new_n873_})
2'b00 : new_n2104_ = 1'b1;
default : new_n2104_ = 1'b0;
endcase
casez ({new_n396_, new_n584_})
2'b00 : new_n2105_ = 1'b1;
default : new_n2105_ = 1'b0;
endcase
casez ({new_n391_, new_n683_})
2'b00 : new_n2106_ = 1'b1;
default : new_n2106_ = 1'b0;
endcase
casez ({new_n442_, new_n717_})
2'b00 : new_n2107_ = 1'b1;
default : new_n2107_ = 1'b0;
endcase
casez ({new_n145_, new_n422_})
2'b00 : new_n2108_ = 1'b1;
default : new_n2108_ = 1'b0;
endcase
casez ({new_n132_, new_n239_})
2'b00 : new_n2109_ = 1'b1;
default : new_n2109_ = 1'b0;
endcase
casez ({new_n109_, new_n799_})
2'b01 : new_n2110_ = 1'b1;
default : new_n2110_ = 1'b0;
endcase
casez ({new_n79_, new_n799_})
2'b01 : new_n2111_ = 1'b1;
default : new_n2111_ = 1'b0;
endcase
casez ({new_n120_, new_n526_})
2'b11 : new_n2112_ = 1'b1;
default : new_n2112_ = 1'b0;
endcase
casez ({x[0], new_n527_})
2'b11 : new_n2113_ = 1'b1;
default : new_n2113_ = 1'b0;
endcase
casez ({new_n91_, new_n542_})
2'b11 : new_n2114_ = 1'b1;
default : new_n2114_ = 1'b0;
endcase
casez ({new_n79_, new_n557_})
2'b11 : new_n2115_ = 1'b1;
default : new_n2115_ = 1'b0;
endcase
casez ({new_n92_, new_n289_})
2'b11 : new_n2116_ = 1'b1;
default : new_n2116_ = 1'b0;
endcase
casez ({u[1], new_n290_})
2'b01 : new_n2117_ = 1'b1;
default : new_n2117_ = 1'b0;
endcase
casez ({new_n83_, new_n292_})
2'b11 : new_n2118_ = 1'b1;
default : new_n2118_ = 1'b0;
endcase
casez ({u[0], new_n295_})
2'b11 : new_n2119_ = 1'b1;
default : new_n2119_ = 1'b0;
endcase
casez ({x[0], new_n295_})
2'b11 : new_n2120_ = 1'b1;
default : new_n2120_ = 1'b0;
endcase
casez ({new_n89_, new_n583_})
2'b11 : new_n2121_ = 1'b1;
default : new_n2121_ = 1'b0;
endcase
casez ({new_n95_, new_n308_})
2'b11 : new_n2122_ = 1'b1;
default : new_n2122_ = 1'b0;
endcase
casez ({new_n77_, new_n308_})
2'b01 : new_n2123_ = 1'b1;
default : new_n2123_ = 1'b0;
endcase
casez ({new_n186_, new_n309_})
2'b11 : new_n2124_ = 1'b1;
default : new_n2124_ = 1'b0;
endcase
casez ({u[0], new_n310_})
2'b11 : new_n2125_ = 1'b1;
default : new_n2125_ = 1'b0;
endcase
casez ({new_n88_, new_n181_})
2'b10 : new_n2126_ = 1'b1;
default : new_n2126_ = 1'b0;
endcase
casez ({v[1], new_n185_})
2'b11 : new_n2127_ = 1'b1;
default : new_n2127_ = 1'b0;
endcase
casez ({new_n148_, new_n186_})
2'b11 : new_n2128_ = 1'b1;
default : new_n2128_ = 1'b0;
endcase
casez ({u[1], new_n330_})
2'b11 : new_n2129_ = 1'b1;
default : new_n2129_ = 1'b0;
endcase
casez ({x[2], new_n330_})
2'b11 : new_n2130_ = 1'b1;
default : new_n2130_ = 1'b0;
endcase
casez ({u[0], new_n335_})
2'b11 : new_n2131_ = 1'b1;
default : new_n2131_ = 1'b0;
endcase
casez ({new_n89_, new_n345_})
2'b11 : new_n2132_ = 1'b1;
default : new_n2132_ = 1'b0;
endcase
casez ({new_n88_, new_n345_})
2'b11 : new_n2133_ = 1'b1;
default : new_n2133_ = 1'b0;
endcase
casez ({u[0], new_n345_})
2'b11 : new_n2134_ = 1'b1;
default : new_n2134_ = 1'b0;
endcase
casez ({new_n88_, new_n352_})
2'b11 : new_n2135_ = 1'b1;
default : new_n2135_ = 1'b0;
endcase
casez ({new_n103_, new_n353_})
2'b11 : new_n2136_ = 1'b1;
default : new_n2136_ = 1'b0;
endcase
casez ({u[0], new_n366_})
2'b01 : new_n2137_ = 1'b1;
default : new_n2137_ = 1'b0;
endcase
casez ({u[1], new_n377_})
2'b11 : new_n2138_ = 1'b1;
default : new_n2138_ = 1'b0;
endcase
casez ({new_n103_, new_n378_})
2'b11 : new_n2139_ = 1'b1;
default : new_n2139_ = 1'b0;
endcase
casez ({new_n88_, new_n382_})
2'b11 : new_n2140_ = 1'b1;
default : new_n2140_ = 1'b0;
endcase
casez ({new_n103_, new_n387_})
2'b11 : new_n2141_ = 1'b1;
default : new_n2141_ = 1'b0;
endcase
casez ({new_n104_, new_n389_})
2'b11 : new_n2142_ = 1'b1;
default : new_n2142_ = 1'b0;
endcase
casez ({y[0], new_n397_})
2'b01 : new_n2143_ = 1'b1;
default : new_n2143_ = 1'b0;
endcase
casez ({new_n215_, new_n398_})
2'b11 : new_n2144_ = 1'b1;
default : new_n2144_ = 1'b0;
endcase
casez ({x[0], new_n404_})
2'b01 : new_n2145_ = 1'b1;
default : new_n2145_ = 1'b0;
endcase
casez ({new_n101_, new_n405_})
2'b11 : new_n2146_ = 1'b1;
default : new_n2146_ = 1'b0;
endcase
casez ({new_n89_, new_n407_})
2'b11 : new_n2147_ = 1'b1;
default : new_n2147_ = 1'b0;
endcase
casez ({new_n150_, new_n418_})
2'b10 : new_n2148_ = 1'b1;
default : new_n2148_ = 1'b0;
endcase
casez ({new_n116_, new_n442_})
2'b11 : new_n2149_ = 1'b1;
default : new_n2149_ = 1'b0;
endcase
casez ({new_n79_, new_n449_})
2'b01 : new_n2150_ = 1'b1;
default : new_n2150_ = 1'b0;
endcase
casez ({x[0], new_n451_})
2'b11 : new_n2151_ = 1'b1;
default : new_n2151_ = 1'b0;
endcase
casez ({new_n79_, new_n457_})
2'b11 : new_n2152_ = 1'b1;
default : new_n2152_ = 1'b0;
endcase
casez ({new_n118_, new_n134_})
2'b11 : new_n2153_ = 1'b1;
default : new_n2153_ = 1'b0;
endcase
casez ({v[1], new_n252_})
2'b00 : new_n2154_ = 1'b1;
default : new_n2154_ = 1'b0;
endcase
casez ({new_n115_, new_n157_})
2'b11 : new_n2155_ = 1'b1;
default : new_n2155_ = 1'b0;
endcase
casez ({x[0], new_n157_})
2'b11 : new_n2156_ = 1'b1;
default : new_n2156_ = 1'b0;
endcase
casez ({new_n83_, new_n265_})
2'b11 : new_n2157_ = 1'b1;
default : new_n2157_ = 1'b0;
endcase
casez ({x[0], new_n175_})
2'b11 : new_n2158_ = 1'b1;
default : new_n2158_ = 1'b0;
endcase
casez ({new_n83_, new_n179_})
2'b11 : new_n2159_ = 1'b1;
default : new_n2159_ = 1'b0;
endcase
casez ({new_n84_, new_n323_})
2'b11 : new_n2160_ = 1'b1;
default : new_n2160_ = 1'b0;
endcase
casez ({new_n84_, new_n134_})
2'b11 : new_n2161_ = 1'b1;
default : new_n2161_ = 1'b0;
endcase
casez ({new_n236_, new_n283_})
2'b00 : new_n2162_ = 1'b1;
default : new_n2162_ = 1'b0;
endcase
casez ({new_n270_, new_n289_})
2'b00 : new_n2163_ = 1'b1;
default : new_n2163_ = 1'b0;
endcase
casez ({new_n269_, new_n311_})
2'b00 : new_n2164_ = 1'b1;
default : new_n2164_ = 1'b0;
endcase
casez ({new_n265_, new_n379_})
2'b00 : new_n2165_ = 1'b1;
default : new_n2165_ = 1'b0;
endcase
casez ({new_n253_, new_n416_})
2'b00 : new_n2166_ = 1'b1;
default : new_n2166_ = 1'b0;
endcase
casez ({new_n5451_, new_n791_, new_n1909_})
3'b1?? : new_n2167_ = 1'b1;
3'b?11 : new_n2167_ = 1'b1;
default : new_n2167_ = 1'b0;
endcase
casez ({new_n250_, new_n649_, new_n472_, new_n771_})
4'b11?? : new_n2168_ = 1'b1;
4'b??11 : new_n2168_ = 1'b1;
default : new_n2168_ = 1'b0;
endcase
casez ({new_n5436_, new_n274_, new_n1149_})
3'b1?? : new_n2169_ = 1'b1;
3'b?11 : new_n2169_ = 1'b1;
default : new_n2169_ = 1'b0;
endcase
casez ({new_n260_, new_n725_, new_n263_, new_n1151_})
4'b11?? : new_n2170_ = 1'b1;
4'b??11 : new_n2170_ = 1'b1;
default : new_n2170_ = 1'b0;
endcase
casez ({new_n162_, new_n907_, new_n216_, new_n1157_})
4'b11?? : new_n2171_ = 1'b1;
4'b??11 : new_n2171_ = 1'b1;
default : new_n2171_ = 1'b0;
endcase
casez ({new_n210_, new_n1499_, new_n350_, new_n1954_})
4'b11?? : new_n2172_ = 1'b1;
4'b??11 : new_n2172_ = 1'b1;
default : new_n2172_ = 1'b0;
endcase
casez ({new_n289_, new_n501_, new_n324_, new_n368_})
4'b11?? : new_n2173_ = 1'b1;
4'b??11 : new_n2173_ = 1'b1;
default : new_n2173_ = 1'b0;
endcase
casez ({new_n437_, new_n1591_, new_n623_, new_n1962_})
4'b11?? : new_n2174_ = 1'b1;
4'b??11 : new_n2174_ = 1'b1;
default : new_n2174_ = 1'b0;
endcase
casez ({new_n149_, new_n269_, new_n270_, new_n793_})
4'b11?? : new_n2175_ = 1'b1;
4'b??11 : new_n2175_ = 1'b1;
default : new_n2175_ = 1'b0;
endcase
casez ({new_n138_, new_n510_, new_n347_, new_n368_})
4'b11?? : new_n2176_ = 1'b1;
4'b??11 : new_n2176_ = 1'b1;
default : new_n2176_ = 1'b0;
endcase
casez ({new_n424_, new_n479_, new_n744_, new_n1181_})
4'b11?? : new_n2177_ = 1'b1;
4'b??11 : new_n2177_ = 1'b1;
default : new_n2177_ = 1'b0;
endcase
casez ({new_n174_, new_n1374_, new_n405_, new_n2012_})
4'b11?? : new_n2178_ = 1'b1;
4'b??10 : new_n2178_ = 1'b1;
default : new_n2178_ = 1'b0;
endcase
casez ({new_n347_, new_n1187_})
2'b01 : new_n2179_ = 1'b1;
default : new_n2179_ = 1'b0;
endcase
casez ({new_n140_, new_n646_, new_n5431_})
3'b11? : new_n2180_ = 1'b1;
3'b??1 : new_n2180_ = 1'b1;
default : new_n2180_ = 1'b0;
endcase
casez ({new_n179_, new_n2039_, new_n229_, new_n945_})
4'b10?? : new_n2181_ = 1'b1;
4'b??11 : new_n2181_ = 1'b1;
default : new_n2181_ = 1'b0;
endcase
casez ({new_n373_, new_n552_, new_n414_, new_n807_})
4'b11?? : new_n2182_ = 1'b1;
4'b??11 : new_n2182_ = 1'b1;
default : new_n2182_ = 1'b0;
endcase
casez ({new_n271_, new_n1281_, new_n603_, new_n2048_})
4'b11?? : new_n2183_ = 1'b1;
4'b??10 : new_n2183_ = 1'b1;
default : new_n2183_ = 1'b0;
endcase
casez ({new_n5446_, new_n508_, new_n1201_})
3'b1?? : new_n2184_ = 1'b1;
3'b?11 : new_n2184_ = 1'b1;
default : new_n2184_ = 1'b0;
endcase
casez ({new_n142_, new_n678_, new_n210_, new_n808_})
4'b11?? : new_n2185_ = 1'b1;
4'b??11 : new_n2185_ = 1'b1;
default : new_n2185_ = 1'b0;
endcase
casez ({new_n142_, new_n1204_, new_n158_, new_n902_})
4'b11?? : new_n2186_ = 1'b1;
4'b??11 : new_n2186_ = 1'b1;
default : new_n2186_ = 1'b0;
endcase
casez ({new_n183_, new_n710_, new_n216_, new_n809_})
4'b11?? : new_n2187_ = 1'b1;
4'b??11 : new_n2187_ = 1'b1;
default : new_n2187_ = 1'b0;
endcase
casez ({new_n986_, new_n1207_})
2'b00 : new_n2188_ = 1'b1;
default : new_n2188_ = 1'b0;
endcase
casez ({new_n129_, new_n1859_, new_n381_, new_n2076_})
4'b11?? : new_n2189_ = 1'b1;
4'b??10 : new_n2189_ = 1'b1;
default : new_n2189_ = 1'b0;
endcase
casez ({new_n368_, new_n2079_, new_n433_, new_n506_})
4'b10?? : new_n2190_ = 1'b1;
4'b??11 : new_n2190_ = 1'b1;
default : new_n2190_ = 1'b0;
endcase
casez ({new_n150_, new_n809_, new_n305_, new_n1208_})
4'b11?? : new_n2191_ = 1'b1;
4'b??11 : new_n2191_ = 1'b1;
default : new_n2191_ = 1'b0;
endcase
casez ({new_n118_, new_n1209_, new_n267_, new_n853_})
4'b11?? : new_n2192_ = 1'b1;
4'b??11 : new_n2192_ = 1'b1;
default : new_n2192_ = 1'b0;
endcase
casez ({new_n86_, new_n464_, new_n115_, new_n1211_})
4'b11?? : new_n2193_ = 1'b1;
4'b??11 : new_n2193_ = 1'b1;
default : new_n2193_ = 1'b0;
endcase
casez ({new_n601_, new_n1211_})
2'b00 : new_n2194_ = 1'b1;
default : new_n2194_ = 1'b0;
endcase
casez ({new_n249_, new_n813_, new_n281_, new_n464_})
4'b11?? : new_n2195_ = 1'b1;
4'b??11 : new_n2195_ = 1'b1;
default : new_n2195_ = 1'b0;
endcase
casez ({new_n216_, new_n611_, new_n263_, new_n1212_})
4'b11?? : new_n2196_ = 1'b1;
4'b??11 : new_n2196_ = 1'b1;
default : new_n2196_ = 1'b0;
endcase
casez ({new_n241_, new_n725_, new_n278_, new_n814_})
4'b11?? : new_n2197_ = 1'b1;
4'b??11 : new_n2197_ = 1'b1;
default : new_n2197_ = 1'b0;
endcase
casez ({new_n300_, new_n814_, new_n317_, new_n649_})
4'b11?? : new_n2198_ = 1'b1;
4'b??11 : new_n2198_ = 1'b1;
default : new_n2198_ = 1'b0;
endcase
casez ({new_n5452_, new_n250_, new_n1214_})
3'b1?? : new_n2199_ = 1'b1;
3'b?11 : new_n2199_ = 1'b1;
default : new_n2199_ = 1'b0;
endcase
casez ({new_n835_, new_n1215_})
2'b00 : new_n2200_ = 1'b1;
default : new_n2200_ = 1'b0;
endcase
casez ({new_n93_, new_n2112_, new_n213_, new_n859_})
4'b11?? : new_n2201_ = 1'b1;
4'b??11 : new_n2201_ = 1'b1;
default : new_n2201_ = 1'b0;
endcase
casez ({new_n104_, new_n1217_, new_n239_, new_n506_})
4'b11?? : new_n2202_ = 1'b1;
4'b??11 : new_n2202_ = 1'b1;
default : new_n2202_ = 1'b0;
endcase
casez ({new_n151_, new_n1217_, new_n284_, new_n808_})
4'b11?? : new_n2203_ = 1'b1;
4'b??11 : new_n2203_ = 1'b1;
default : new_n2203_ = 1'b0;
endcase
casez ({new_n278_, new_n1555_, new_n284_, new_n2115_})
4'b11?? : new_n2204_ = 1'b1;
4'b??11 : new_n2204_ = 1'b1;
default : new_n2204_ = 1'b0;
endcase
casez ({new_n86_, new_n482_, new_n243_, new_n1219_})
4'b11?? : new_n2205_ = 1'b1;
4'b??11 : new_n2205_ = 1'b1;
default : new_n2205_ = 1'b0;
endcase
casez ({new_n113_, new_n1223_, new_n279_, new_n2120_})
4'b11?? : new_n2206_ = 1'b1;
4'b??11 : new_n2206_ = 1'b1;
default : new_n2206_ = 1'b0;
endcase
casez ({new_n84_, new_n2123_, new_n172_, new_n899_})
4'b11?? : new_n2207_ = 1'b1;
4'b??11 : new_n2207_ = 1'b1;
default : new_n2207_ = 1'b0;
endcase
casez ({new_n239_, new_n2127_, new_n306_, new_n1468_})
4'b11?? : new_n2208_ = 1'b1;
4'b??11 : new_n2208_ = 1'b1;
default : new_n2208_ = 1'b0;
endcase
casez ({new_n309_, new_n2129_, new_n5443_})
3'b11? : new_n2209_ = 1'b1;
3'b??1 : new_n2209_ = 1'b1;
default : new_n2209_ = 1'b0;
endcase
casez ({new_n178_, new_n1226_, new_n226_, new_n737_})
4'b11?? : new_n2210_ = 1'b1;
4'b??11 : new_n2210_ = 1'b1;
default : new_n2210_ = 1'b0;
endcase
casez ({new_n127_, new_n1206_, new_n527_, new_n1228_})
4'b11?? : new_n2211_ = 1'b1;
4'b??11 : new_n2211_ = 1'b1;
default : new_n2211_ = 1'b0;
endcase
casez ({new_n305_, new_n981_, new_n433_, new_n2133_})
4'b11?? : new_n2212_ = 1'b1;
4'b??11 : new_n2212_ = 1'b1;
default : new_n2212_ = 1'b0;
endcase
casez ({new_n167_, new_n833_, new_n246_, new_n2134_})
4'b11?? : new_n2213_ = 1'b1;
4'b??11 : new_n2213_ = 1'b1;
default : new_n2213_ = 1'b0;
endcase
casez ({new_n118_, new_n2135_, new_n167_, new_n838_})
4'b11?? : new_n2214_ = 1'b1;
4'b??11 : new_n2214_ = 1'b1;
default : new_n2214_ = 1'b0;
endcase
casez ({new_n164_, new_n1823_, new_n493_, new_n2142_})
4'b11?? : new_n2215_ = 1'b1;
4'b??11 : new_n2215_ = 1'b1;
default : new_n2215_ = 1'b0;
endcase
casez ({new_n201_, new_n832_, new_n224_, new_n828_})
4'b11?? : new_n2216_ = 1'b1;
4'b??11 : new_n2216_ = 1'b1;
default : new_n2216_ = 1'b0;
endcase
casez ({new_n167_, new_n1284_, new_n438_, new_n2147_})
4'b11?? : new_n2217_ = 1'b1;
4'b??11 : new_n2217_ = 1'b1;
default : new_n2217_ = 1'b0;
endcase
casez ({new_n5434_, new_n210_, new_n573_})
3'b1?? : new_n2218_ = 1'b1;
3'b?11 : new_n2218_ = 1'b1;
default : new_n2218_ = 1'b0;
endcase
casez ({new_n800_, new_n842_})
2'b00 : new_n2219_ = 1'b1;
default : new_n2219_ = 1'b0;
endcase
casez ({new_n122_, new_n755_, new_n159_, new_n844_})
4'b11?? : new_n2220_ = 1'b1;
4'b??11 : new_n2220_ = 1'b1;
default : new_n2220_ = 1'b0;
endcase
casez ({new_n160_, new_n852_, new_n187_, new_n647_})
4'b11?? : new_n2221_ = 1'b1;
4'b??11 : new_n2221_ = 1'b1;
default : new_n2221_ = 1'b0;
endcase
casez ({new_n645_, new_n1266_})
2'b00 : new_n2222_ = 1'b1;
default : new_n2222_ = 1'b0;
endcase
casez ({new_n134_, new_n561_, new_n426_, new_n462_})
4'b11?? : new_n2223_ = 1'b1;
4'b??11 : new_n2223_ = 1'b1;
default : new_n2223_ = 1'b0;
endcase
casez ({new_n754_, new_n861_})
2'b00 : new_n2224_ = 1'b1;
default : new_n2224_ = 1'b0;
endcase
casez ({new_n190_, new_n193_, new_n304_, new_n561_})
4'b11?? : new_n2225_ = 1'b1;
4'b??01 : new_n2225_ = 1'b1;
default : new_n2225_ = 1'b0;
endcase
casez ({new_n462_, new_n1268_})
2'b00 : new_n2226_ = 1'b1;
default : new_n2226_ = 1'b0;
endcase
casez ({new_n202_, new_n1271_, new_n230_, new_n513_})
4'b11?? : new_n2227_ = 1'b1;
4'b??11 : new_n2227_ = 1'b1;
default : new_n2227_ = 1'b0;
endcase
casez ({new_n219_, new_n1061_, new_n241_, new_n1286_})
4'b11?? : new_n2228_ = 1'b1;
4'b??11 : new_n2228_ = 1'b1;
default : new_n2228_ = 1'b0;
endcase
casez ({new_n5448_, new_n538_, new_n1289_})
3'b1?? : new_n2229_ = 1'b1;
3'b?11 : new_n2229_ = 1'b1;
default : new_n2229_ = 1'b0;
endcase
casez ({new_n161_, new_n1291_, new_n305_, new_n647_})
4'b11?? : new_n2230_ = 1'b1;
4'b??11 : new_n2230_ = 1'b1;
default : new_n2230_ = 1'b0;
endcase
casez ({new_n222_, new_n1297_, new_n267_, new_n983_})
4'b11?? : new_n2231_ = 1'b1;
4'b??11 : new_n2231_ = 1'b1;
default : new_n2231_ = 1'b0;
endcase
casez ({new_n171_, new_n567_, new_n174_, new_n514_})
4'b11?? : new_n2232_ = 1'b1;
4'b??11 : new_n2232_ = 1'b1;
default : new_n2232_ = 1'b0;
endcase
casez ({new_n214_, new_n1308_, new_n287_, new_n611_})
4'b11?? : new_n2233_ = 1'b1;
4'b??11 : new_n2233_ = 1'b1;
default : new_n2233_ = 1'b0;
endcase
casez ({new_n5455_, new_n729_, new_n1315_})
3'b1?? : new_n2234_ = 1'b1;
3'b?11 : new_n2234_ = 1'b1;
default : new_n2234_ = 1'b0;
endcase
casez ({new_n113_, new_n662_, new_n252_, new_n1317_})
4'b11?? : new_n2235_ = 1'b1;
4'b??01 : new_n2235_ = 1'b1;
default : new_n2235_ = 1'b0;
endcase
casez ({new_n148_, new_n907_, new_n151_, new_n1318_})
4'b11?? : new_n2236_ = 1'b1;
4'b??11 : new_n2236_ = 1'b1;
default : new_n2236_ = 1'b0;
endcase
casez ({new_n791_, new_n1321_})
2'b00 : new_n2237_ = 1'b1;
default : new_n2237_ = 1'b0;
endcase
casez ({new_n104_, new_n575_, new_n120_, new_n277_})
4'b11?? : new_n2238_ = 1'b1;
4'b??11 : new_n2238_ = 1'b1;
default : new_n2238_ = 1'b0;
endcase
casez ({new_n290_, new_n1331_, new_n381_, new_n1028_})
4'b11?? : new_n2239_ = 1'b1;
4'b??11 : new_n2239_ = 1'b1;
default : new_n2239_ = 1'b0;
endcase
casez ({new_n138_, new_n610_, new_n633_, new_n1335_})
4'b11?? : new_n2240_ = 1'b1;
4'b??11 : new_n2240_ = 1'b1;
default : new_n2240_ = 1'b0;
endcase
casez ({new_n696_, new_n1339_})
2'b00 : new_n2241_ = 1'b1;
default : new_n2241_ = 1'b0;
endcase
casez ({new_n168_, new_n1342_, new_n170_, new_n1104_})
4'b11?? : new_n2242_ = 1'b1;
4'b??11 : new_n2242_ = 1'b1;
default : new_n2242_ = 1'b0;
endcase
casez ({new_n544_, new_n1353_})
2'b00 : new_n2243_ = 1'b1;
default : new_n2243_ = 1'b0;
endcase
casez ({new_n245_, new_n897_})
2'b00 : new_n2244_ = 1'b1;
default : new_n2244_ = 1'b0;
endcase
casez ({new_n152_, new_n898_, new_n270_, new_n538_})
4'b11?? : new_n2245_ = 1'b1;
4'b??11 : new_n2245_ = 1'b1;
default : new_n2245_ = 1'b0;
endcase
casez ({new_n274_, new_n1360_, new_n462_, new_n794_})
4'b11?? : new_n2246_ = 1'b1;
4'b??11 : new_n2246_ = 1'b1;
default : new_n2246_ = 1'b0;
endcase
casez ({new_n155_, new_n900_, new_n214_, new_n723_})
4'b11?? : new_n2247_ = 1'b1;
4'b??11 : new_n2247_ = 1'b1;
default : new_n2247_ = 1'b0;
endcase
casez ({new_n189_, new_n720_, new_n213_, new_n901_})
4'b10?? : new_n2248_ = 1'b1;
4'b??11 : new_n2248_ = 1'b1;
default : new_n2248_ = 1'b0;
endcase
casez ({new_n240_, new_n613_, new_n381_, new_n1367_})
4'b11?? : new_n2249_ = 1'b1;
4'b??11 : new_n2249_ = 1'b1;
default : new_n2249_ = 1'b0;
endcase
casez ({new_n91_, new_n699_, new_n385_, new_n902_})
4'b11?? : new_n2250_ = 1'b1;
4'b??11 : new_n2250_ = 1'b1;
default : new_n2250_ = 1'b0;
endcase
casez ({new_n182_, new_n1372_, new_n979_, new_n1126_})
4'b11?? : new_n2251_ = 1'b1;
4'b??11 : new_n2251_ = 1'b1;
default : new_n2251_ = 1'b0;
endcase
casez ({new_n142_, new_n904_, new_n164_, new_n295_})
4'b11?? : new_n2252_ = 1'b1;
4'b??11 : new_n2252_ = 1'b1;
default : new_n2252_ = 1'b0;
endcase
casez ({new_n442_, new_n906_, new_n612_, new_n709_})
4'b11?? : new_n2253_ = 1'b1;
4'b??10 : new_n2253_ = 1'b1;
default : new_n2253_ = 1'b0;
endcase
casez ({new_n1218_, new_n1384_})
2'b00 : new_n2254_ = 1'b1;
default : new_n2254_ = 1'b0;
endcase
casez ({new_n89_, new_n909_, new_n222_, new_n699_})
4'b11?? : new_n2255_ = 1'b1;
4'b??11 : new_n2255_ = 1'b1;
default : new_n2255_ = 1'b0;
endcase
casez ({new_n149_, new_n368_, new_n174_, new_n610_})
4'b11?? : new_n2256_ = 1'b1;
4'b??11 : new_n2256_ = 1'b1;
default : new_n2256_ = 1'b0;
endcase
casez ({new_n237_, new_n695_, new_n387_, new_n1388_})
4'b11?? : new_n2257_ = 1'b1;
4'b??11 : new_n2257_ = 1'b1;
default : new_n2257_ = 1'b0;
endcase
casez ({new_n144_, new_n463_, new_n355_, new_n1412_})
4'b11?? : new_n2258_ = 1'b1;
4'b??10 : new_n2258_ = 1'b1;
default : new_n2258_ = 1'b0;
endcase
casez ({new_n938_, new_n1433_})
2'b01 : new_n2259_ = 1'b1;
default : new_n2259_ = 1'b0;
endcase
casez ({new_n256_, new_n940_})
2'b00 : new_n2260_ = 1'b1;
default : new_n2260_ = 1'b0;
endcase
casez ({new_n624_, new_n941_})
2'b00 : new_n2261_ = 1'b1;
default : new_n2261_ = 1'b0;
endcase
casez ({new_n177_, new_n1457_, new_n4663_})
3'b11? : new_n2262_ = 1'b1;
3'b??1 : new_n2262_ = 1'b1;
default : new_n2262_ = 1'b0;
endcase
casez ({new_n275_, new_n1458_, new_n284_, new_n1056_})
4'b11?? : new_n2263_ = 1'b1;
4'b??11 : new_n2263_ = 1'b1;
default : new_n2263_ = 1'b0;
endcase
casez ({new_n167_, new_n1357_, new_n264_, new_n1458_})
4'b11?? : new_n2264_ = 1'b1;
4'b??11 : new_n2264_ = 1'b1;
default : new_n2264_ = 1'b0;
endcase
casez ({new_n905_, new_n1460_})
2'b00 : new_n2265_ = 1'b1;
default : new_n2265_ = 1'b0;
endcase
casez ({new_n155_, new_n1460_, new_n464_, new_n628_})
4'b11?? : new_n2266_ = 1'b1;
4'b??10 : new_n2266_ = 1'b1;
default : new_n2266_ = 1'b0;
endcase
casez ({new_n477_, new_n1461_})
2'b00 : new_n2267_ = 1'b1;
default : new_n2267_ = 1'b0;
endcase
casez ({new_n90_, new_n624_, new_n205_, new_n1468_})
4'b11?? : new_n2268_ = 1'b1;
4'b??11 : new_n2268_ = 1'b1;
default : new_n2268_ = 1'b0;
endcase
casez ({new_n164_, new_n948_, new_n322_, new_n416_})
4'b11?? : new_n2269_ = 1'b1;
4'b??11 : new_n2269_ = 1'b1;
default : new_n2269_ = 1'b0;
endcase
casez ({new_n139_, new_n1471_, new_n175_, new_n540_})
4'b11?? : new_n2270_ = 1'b1;
4'b??11 : new_n2270_ = 1'b1;
default : new_n2270_ = 1'b0;
endcase
casez ({new_n283_, new_n1405_, new_n469_, new_n1473_})
4'b10?? : new_n2271_ = 1'b1;
4'b??11 : new_n2271_ = 1'b1;
default : new_n2271_ = 1'b0;
endcase
casez ({new_n183_, new_n1477_, new_n355_, new_n1395_})
4'b11?? : new_n2272_ = 1'b1;
4'b??11 : new_n2272_ = 1'b1;
default : new_n2272_ = 1'b0;
endcase
casez ({new_n698_, new_n954_})
2'b00 : new_n2273_ = 1'b1;
default : new_n2273_ = 1'b0;
endcase
casez ({new_n184_, new_n1060_, new_n266_, new_n1479_})
4'b11?? : new_n2274_ = 1'b1;
4'b??11 : new_n2274_ = 1'b1;
default : new_n2274_ = 1'b0;
endcase
casez ({new_n168_, new_n1484_, new_n388_, new_n1065_})
4'b11?? : new_n2275_ = 1'b1;
4'b??11 : new_n2275_ = 1'b1;
default : new_n2275_ = 1'b0;
endcase
casez ({new_n190_, new_n613_, new_n246_, new_n639_})
4'b11?? : new_n2276_ = 1'b1;
4'b??11 : new_n2276_ = 1'b1;
default : new_n2276_ = 1'b0;
endcase
casez ({new_n1203_, new_n1487_})
2'b00 : new_n2277_ = 1'b1;
default : new_n2277_ = 1'b0;
endcase
casez ({new_n187_, new_n1491_, new_n214_, new_n1375_})
4'b11?? : new_n2278_ = 1'b1;
4'b??11 : new_n2278_ = 1'b1;
default : new_n2278_ = 1'b0;
endcase
casez ({new_n159_, new_n643_, new_n427_, new_n506_})
4'b11?? : new_n2279_ = 1'b1;
4'b??11 : new_n2279_ = 1'b1;
default : new_n2279_ = 1'b0;
endcase
casez ({new_n163_, new_n1494_, new_n384_, new_n615_})
4'b11?? : new_n2280_ = 1'b1;
4'b??10 : new_n2280_ = 1'b1;
default : new_n2280_ = 1'b0;
endcase
casez ({new_n5441_, new_n262_, new_n1495_})
3'b1?? : new_n2281_ = 1'b1;
3'b?11 : new_n2281_ = 1'b1;
default : new_n2281_ = 1'b0;
endcase
casez ({new_n1057_, new_n1495_})
2'b00 : new_n2282_ = 1'b1;
default : new_n2282_ = 1'b0;
endcase
casez ({new_n133_, new_n1496_, new_n251_, new_n722_})
4'b11?? : new_n2283_ = 1'b1;
4'b??11 : new_n2283_ = 1'b1;
default : new_n2283_ = 1'b0;
endcase
casez ({new_n85_, new_n757_, new_n90_, new_n1497_})
4'b11?? : new_n2284_ = 1'b1;
4'b??11 : new_n2284_ = 1'b1;
default : new_n2284_ = 1'b0;
endcase
casez ({new_n155_, new_n644_, new_n188_, new_n286_})
4'b11?? : new_n2285_ = 1'b1;
4'b??11 : new_n2285_ = 1'b1;
default : new_n2285_ = 1'b0;
endcase
casez ({new_n218_, new_n1500_, new_n669_, new_n1228_})
4'b11?? : new_n2286_ = 1'b1;
4'b??11 : new_n2286_ = 1'b1;
default : new_n2286_ = 1'b0;
endcase
casez ({new_n494_, new_n973_})
2'b00 : new_n2287_ = 1'b1;
default : new_n2287_ = 1'b0;
endcase
casez ({new_n263_, new_n1505_, new_n346_, new_n1070_})
4'b11?? : new_n2288_ = 1'b1;
4'b??11 : new_n2288_ = 1'b1;
default : new_n2288_ = 1'b0;
endcase
casez ({new_n122_, new_n977_, new_n149_, new_n897_})
4'b11?? : new_n2289_ = 1'b1;
4'b??11 : new_n2289_ = 1'b1;
default : new_n2289_ = 1'b0;
endcase
casez ({new_n89_, new_n978_, new_n137_, new_n939_})
4'b11?? : new_n2290_ = 1'b1;
4'b??11 : new_n2290_ = 1'b1;
default : new_n2290_ = 1'b0;
endcase
casez ({new_n202_, new_n996_, new_n254_, new_n847_})
4'b11?? : new_n2291_ = 1'b1;
4'b??11 : new_n2291_ = 1'b1;
default : new_n2291_ = 1'b0;
endcase
casez ({new_n572_, new_n1567_})
2'b00 : new_n2292_ = 1'b1;
default : new_n2292_ = 1'b0;
endcase
casez ({new_n1060_, new_n1571_})
2'b00 : new_n2293_ = 1'b1;
default : new_n2293_ = 1'b0;
endcase
casez ({new_n222_, new_n1008_, new_n5450_})
3'b11? : new_n2294_ = 1'b1;
3'b??1 : new_n2294_ = 1'b1;
default : new_n2294_ = 1'b0;
endcase
casez ({new_n5447_, new_n311_, new_n426_})
3'b1?? : new_n2295_ = 1'b1;
3'b?11 : new_n2295_ = 1'b1;
default : new_n2295_ = 1'b0;
endcase
casez ({new_n161_, new_n464_, new_n202_, new_n675_})
4'b11?? : new_n2296_ = 1'b1;
4'b??11 : new_n2296_ = 1'b1;
default : new_n2296_ = 1'b0;
endcase
casez ({new_n172_, new_n1586_, new_n179_, new_n726_})
4'b11?? : new_n2297_ = 1'b1;
4'b??11 : new_n2297_ = 1'b1;
default : new_n2297_ = 1'b0;
endcase
casez ({new_n168_, new_n639_, new_n307_, new_n677_})
4'b11?? : new_n2298_ = 1'b1;
4'b??11 : new_n2298_ = 1'b1;
default : new_n2298_ = 1'b0;
endcase
casez ({new_n506_, new_n1012_})
2'b00 : new_n2299_ = 1'b1;
default : new_n2299_ = 1'b0;
endcase
casez ({new_n222_, new_n1597_, new_n344_, new_n661_})
4'b11?? : new_n2300_ = 1'b1;
4'b??11 : new_n2300_ = 1'b1;
default : new_n2300_ = 1'b0;
endcase
casez ({new_n815_, new_n1605_})
2'b00 : new_n2301_ = 1'b1;
default : new_n2301_ = 1'b0;
endcase
casez ({new_n561_, new_n1608_})
2'b00 : new_n2302_ = 1'b1;
default : new_n2302_ = 1'b0;
endcase
casez ({new_n5455_, new_n353_, new_n1610_})
3'b1?? : new_n2303_ = 1'b1;
3'b?11 : new_n2303_ = 1'b1;
default : new_n2303_ = 1'b0;
endcase
casez ({new_n726_, new_n1617_})
2'b00 : new_n2304_ = 1'b1;
default : new_n2304_ = 1'b0;
endcase
casez ({new_n4660_, new_n412_, new_n815_})
3'b1?? : new_n2305_ = 1'b1;
3'b?11 : new_n2305_ = 1'b1;
default : new_n2305_ = 1'b0;
endcase
casez ({u[1], new_n625_, new_n336_, new_n697_})
4'b01?? : new_n2306_ = 1'b1;
4'b??11 : new_n2306_ = 1'b1;
default : new_n2306_ = 1'b0;
endcase
casez ({new_n201_, new_n710_, new_n269_, new_n552_})
4'b11?? : new_n2307_ = 1'b1;
4'b??11 : new_n2307_ = 1'b1;
default : new_n2307_ = 1'b0;
endcase
casez ({new_n192_, new_n942_, new_n221_, new_n1057_})
4'b11?? : new_n2308_ = 1'b1;
4'b??11 : new_n2308_ = 1'b1;
default : new_n2308_ = 1'b0;
endcase
casez ({new_n611_, new_n1058_})
2'b00 : new_n2309_ = 1'b1;
default : new_n2309_ = 1'b0;
endcase
casez ({new_n131_, new_n1058_, new_n342_, new_n699_})
4'b11?? : new_n2310_ = 1'b1;
4'b??11 : new_n2310_ = 1'b1;
default : new_n2310_ = 1'b0;
endcase
casez ({new_n131_, new_n681_, new_n241_, new_n1713_})
4'b11?? : new_n2311_ = 1'b1;
4'b??11 : new_n2311_ = 1'b1;
default : new_n2311_ = 1'b0;
endcase
casez ({new_n1319_, new_n1720_})
2'b00 : new_n2312_ = 1'b1;
default : new_n2312_ = 1'b0;
endcase
casez ({new_n172_, new_n1112_, new_n267_, new_n1720_})
4'b11?? : new_n2313_ = 1'b1;
4'b??11 : new_n2313_ = 1'b1;
default : new_n2313_ = 1'b0;
endcase
casez ({new_n319_, new_n367_, new_n493_, new_n1064_})
4'b01?? : new_n2314_ = 1'b1;
4'b??11 : new_n2314_ = 1'b1;
default : new_n2314_ = 1'b0;
endcase
casez ({new_n256_, new_n722_, new_n536_, new_n695_})
4'b11?? : new_n2315_ = 1'b1;
4'b??11 : new_n2315_ = 1'b1;
default : new_n2315_ = 1'b0;
endcase
casez ({new_n139_, new_n1067_, new_n216_, new_n724_})
4'b11?? : new_n2316_ = 1'b1;
4'b??11 : new_n2316_ = 1'b1;
default : new_n2316_ = 1'b0;
endcase
casez ({new_n722_, new_n1071_})
2'b00 : new_n2317_ = 1'b1;
default : new_n2317_ = 1'b0;
endcase
casez ({new_n367_, new_n726_})
2'b00 : new_n2318_ = 1'b1;
default : new_n2318_ = 1'b0;
endcase
casez ({new_n267_, new_n1743_, new_n540_, new_n629_})
4'b11?? : new_n2319_ = 1'b1;
4'b??10 : new_n2319_ = 1'b1;
default : new_n2319_ = 1'b0;
endcase
casez ({new_n150_, new_n1219_, new_n5449_})
3'b11? : new_n2320_ = 1'b1;
3'b??1 : new_n2320_ = 1'b1;
default : new_n2320_ = 1'b0;
endcase
casez ({new_n168_, new_n1601_, new_n179_, new_n1754_})
4'b11?? : new_n2321_ = 1'b1;
4'b??11 : new_n2321_ = 1'b1;
default : new_n2321_ = 1'b0;
endcase
casez ({new_n304_, new_n1488_, new_n453_, new_n1809_})
4'b01?? : new_n2322_ = 1'b1;
4'b??10 : new_n2322_ = 1'b1;
default : new_n2322_ = 1'b0;
endcase
casez ({new_n277_, new_n2959_, new_n1817_})
3'b11? : new_n2323_ = 1'b1;
3'b??1 : new_n2323_ = 1'b1;
default : new_n2323_ = 1'b0;
endcase
casez ({new_n1171_, new_n1822_, new_n1224_, new_n1750_})
4'b11?? : new_n2324_ = 1'b1;
4'b??11 : new_n2324_ = 1'b1;
default : new_n2324_ = 1'b0;
endcase
casez ({new_n123_, new_n1828_, new_n1496_, new_n1570_})
4'b11?? : new_n2325_ = 1'b1;
4'b??11 : new_n2325_ = 1'b1;
default : new_n2325_ = 1'b0;
endcase
casez ({new_n699_, new_n1116_})
2'b00 : new_n2326_ = 1'b1;
default : new_n2326_ = 1'b0;
endcase
casez ({new_n218_, new_n726_, new_n285_, new_n1117_})
4'b11?? : new_n2327_ = 1'b1;
4'b??11 : new_n2327_ = 1'b1;
default : new_n2327_ = 1'b0;
endcase
casez ({new_n905_, new_n1117_})
2'b00 : new_n2328_ = 1'b1;
default : new_n2328_ = 1'b0;
endcase
casez ({new_n153_, new_n1066_, new_n199_, new_n1120_})
4'b11?? : new_n2329_ = 1'b1;
4'b??11 : new_n2329_ = 1'b1;
default : new_n2329_ = 1'b0;
endcase
casez ({new_n177_, new_n808_, new_n196_, new_n1842_})
4'b11?? : new_n2330_ = 1'b1;
4'b??11 : new_n2330_ = 1'b1;
default : new_n2330_ = 1'b0;
endcase
casez ({new_n277_, new_n1851_, new_n1220_, new_n1545_})
4'b11?? : new_n2331_ = 1'b1;
4'b??11 : new_n2331_ = 1'b1;
default : new_n2331_ = 1'b0;
endcase
casez ({new_n212_, new_n1068_, new_n214_, new_n1861_})
4'b11?? : new_n2332_ = 1'b1;
4'b??11 : new_n2332_ = 1'b1;
default : new_n2332_ = 1'b0;
endcase
casez ({new_n153_, new_n1713_, new_n356_, new_n1873_})
4'b11?? : new_n2333_ = 1'b1;
4'b??11 : new_n2333_ = 1'b1;
default : new_n2333_ = 1'b0;
endcase
casez ({new_n83_, new_n277_})
2'b11 : new_n2334_ = 1'b1;
default : new_n2334_ = 1'b0;
endcase
casez ({new_n92_, new_n312_})
2'b11 : new_n2335_ = 1'b1;
default : new_n2335_ = 1'b0;
endcase
casez ({new_n79_, new_n416_})
2'b11 : new_n2336_ = 1'b1;
default : new_n2336_ = 1'b0;
endcase
casez ({new_n335_, new_n591_})
2'b00 : new_n2337_ = 1'b1;
default : new_n2337_ = 1'b0;
endcase
casez ({new_n689_, new_n1147_})
2'b00 : new_n2338_ = 1'b1;
default : new_n2338_ = 1'b0;
endcase
casez ({new_n468_, new_n778_})
2'b00 : new_n2339_ = 1'b1;
default : new_n2339_ = 1'b0;
endcase
casez ({new_n219_, new_n258_, new_n394_, new_n1938_})
4'b110? : new_n2340_ = 1'b1;
4'b???1 : new_n2340_ = 1'b1;
default : new_n2340_ = 1'b0;
endcase
casez ({new_n481_, new_n3535_, new_n1967_})
3'b11? : new_n2341_ = 1'b1;
3'b??1 : new_n2341_ = 1'b1;
default : new_n2341_ = 1'b0;
endcase
casez ({new_n299_, new_n2954_, new_n1970_})
3'b11? : new_n2342_ = 1'b1;
3'b??1 : new_n2342_ = 1'b1;
default : new_n2342_ = 1'b0;
endcase
casez ({new_n89_, new_n205_, new_n494_, new_n1972_})
4'b111? : new_n2343_ = 1'b1;
4'b???1 : new_n2343_ = 1'b1;
default : new_n2343_ = 1'b0;
endcase
casez ({new_n204_, new_n219_, new_n222_, new_n1973_})
4'b111? : new_n2344_ = 1'b1;
4'b???1 : new_n2344_ = 1'b1;
default : new_n2344_ = 1'b0;
endcase
casez ({new_n167_, new_n250_, new_n969_, new_n1974_})
4'b110? : new_n2345_ = 1'b1;
4'b???1 : new_n2345_ = 1'b1;
default : new_n2345_ = 1'b0;
endcase
casez ({new_n467_, new_n3478_, new_n1978_})
3'b11? : new_n2346_ = 1'b1;
3'b??1 : new_n2346_ = 1'b1;
default : new_n2346_ = 1'b0;
endcase
casez ({new_n483_, new_n3510_, new_n1979_})
3'b11? : new_n2347_ = 1'b1;
3'b??1 : new_n2347_ = 1'b1;
default : new_n2347_ = 1'b0;
endcase
casez ({new_n314_, new_n2935_, new_n1987_})
3'b11? : new_n2348_ = 1'b1;
3'b??1 : new_n2348_ = 1'b1;
default : new_n2348_ = 1'b0;
endcase
casez ({new_n289_, new_n2947_, new_n1991_})
3'b11? : new_n2349_ = 1'b1;
3'b??1 : new_n2349_ = 1'b1;
default : new_n2349_ = 1'b0;
endcase
casez ({new_n223_, new_n547_, new_n279_, new_n1178_})
4'b11?? : new_n2350_ = 1'b1;
4'b??11 : new_n2350_ = 1'b1;
default : new_n2350_ = 1'b0;
endcase
casez ({new_n265_, new_n3503_, new_n1993_})
3'b11? : new_n2351_ = 1'b1;
3'b??1 : new_n2351_ = 1'b1;
default : new_n2351_ = 1'b0;
endcase
casez ({new_n96_, new_n267_, new_n366_, new_n1996_})
4'b111? : new_n2352_ = 1'b1;
4'b???1 : new_n2352_ = 1'b1;
default : new_n2352_ = 1'b0;
endcase
casez ({y[2], new_n283_, new_n313_, new_n2003_})
4'b011? : new_n2353_ = 1'b1;
4'b???1 : new_n2353_ = 1'b1;
default : new_n2353_ = 1'b0;
endcase
casez ({new_n86_, new_n4624_, new_n2005_})
3'b11? : new_n2354_ = 1'b1;
3'b??1 : new_n2354_ = 1'b1;
default : new_n2354_ = 1'b0;
endcase
casez ({new_n246_, new_n3325_, new_n2011_})
3'b11? : new_n2355_ = 1'b1;
3'b??1 : new_n2355_ = 1'b1;
default : new_n2355_ = 1'b0;
endcase
casez ({new_n320_, new_n3371_, new_n2010_})
3'b01? : new_n2356_ = 1'b1;
3'b??1 : new_n2356_ = 1'b1;
default : new_n2356_ = 1'b0;
endcase
casez ({new_n89_, new_n217_, new_n441_, new_n2015_})
4'b111? : new_n2357_ = 1'b1;
4'b???1 : new_n2357_ = 1'b1;
default : new_n2357_ = 1'b0;
endcase
casez ({new_n716_, new_n4659_, new_n1188_})
3'b11? : new_n2358_ = 1'b1;
3'b??1 : new_n2358_ = 1'b1;
default : new_n2358_ = 1'b0;
endcase
casez ({new_n127_, new_n3452_, new_n2025_})
3'b11? : new_n2359_ = 1'b1;
3'b??1 : new_n2359_ = 1'b1;
default : new_n2359_ = 1'b0;
endcase
casez ({new_n175_, new_n3417_, new_n2031_})
3'b11? : new_n2360_ = 1'b1;
3'b??1 : new_n2360_ = 1'b1;
default : new_n2360_ = 1'b0;
endcase
casez ({new_n95_, new_n150_, new_n251_, new_n1196_})
4'b111? : new_n2361_ = 1'b1;
4'b???1 : new_n2361_ = 1'b1;
default : new_n2361_ = 1'b0;
endcase
casez ({new_n426_, new_n3593_, new_n2037_})
3'b11? : new_n2362_ = 1'b1;
3'b??1 : new_n2362_ = 1'b1;
default : new_n2362_ = 1'b0;
endcase
casez ({new_n591_, new_n803_})
2'b00 : new_n2363_ = 1'b1;
default : new_n2363_ = 1'b0;
endcase
casez ({new_n204_, new_n211_, new_n225_, new_n2045_})
4'b111? : new_n2364_ = 1'b1;
4'b???1 : new_n2364_ = 1'b1;
default : new_n2364_ = 1'b0;
endcase
casez ({v[1], new_n261_, new_n1182_, new_n2056_})
4'b111? : new_n2365_ = 1'b1;
4'b???1 : new_n2365_ = 1'b1;
default : new_n2365_ = 1'b0;
endcase
casez ({x[1], new_n145_, new_n1650_, new_n2070_})
4'b111? : new_n2366_ = 1'b1;
4'b???1 : new_n2366_ = 1'b1;
default : new_n2366_ = 1'b0;
endcase
casez ({new_n95_, new_n207_, new_n449_, new_n2073_})
4'b111? : new_n2367_ = 1'b1;
4'b???1 : new_n2367_ = 1'b1;
default : new_n2367_ = 1'b0;
endcase
casez ({new_n98_, new_n140_, new_n497_, new_n2074_})
4'b111? : new_n2368_ = 1'b1;
4'b???1 : new_n2368_ = 1'b1;
default : new_n2368_ = 1'b0;
endcase
casez ({new_n255_, new_n4590_, new_n2083_})
3'b11? : new_n2369_ = 1'b1;
3'b??1 : new_n2369_ = 1'b1;
default : new_n2369_ = 1'b0;
endcase
casez ({x[2], new_n216_, new_n634_, new_n2084_})
4'b011? : new_n2370_ = 1'b1;
4'b???1 : new_n2370_ = 1'b1;
default : new_n2370_ = 1'b0;
endcase
casez ({new_n372_, new_n3577_, new_n2092_})
3'b11? : new_n2371_ = 1'b1;
3'b??1 : new_n2371_ = 1'b1;
default : new_n2371_ = 1'b0;
endcase
casez ({new_n161_, new_n3334_, new_n2096_})
3'b11? : new_n2372_ = 1'b1;
3'b??1 : new_n2372_ = 1'b1;
default : new_n2372_ = 1'b0;
endcase
casez ({new_n151_, new_n570_, new_n242_, new_n819_})
4'b11?? : new_n2373_ = 1'b1;
4'b??11 : new_n2373_ = 1'b1;
default : new_n2373_ = 1'b0;
endcase
casez ({new_n414_, new_n563_, new_n432_, new_n2123_})
4'b11?? : new_n2374_ = 1'b1;
4'b??11 : new_n2374_ = 1'b1;
default : new_n2374_ = 1'b0;
endcase
casez ({new_n5920_, new_n461_, new_n815_})
3'b1?? : new_n2375_ = 1'b1;
3'b?11 : new_n2375_ = 1'b1;
default : new_n2375_ = 1'b0;
endcase
casez ({new_n166_, new_n640_, new_n194_, new_n2141_})
4'b11?? : new_n2376_ = 1'b1;
4'b??11 : new_n2376_ = 1'b1;
default : new_n2376_ = 1'b0;
endcase
casez ({new_n159_, new_n547_, new_n278_, new_n468_})
4'b11?? : new_n2377_ = 1'b1;
4'b??11 : new_n2377_ = 1'b1;
default : new_n2377_ = 1'b0;
endcase
casez ({new_n103_, new_n547_, new_n178_, new_n518_})
4'b11?? : new_n2378_ = 1'b1;
4'b??11 : new_n2378_ = 1'b1;
default : new_n2378_ = 1'b0;
endcase
casez ({new_n1229_, new_n2162_})
2'b11 : new_n2379_ = 1'b1;
default : new_n2379_ = 1'b0;
endcase
casez ({new_n170_, new_n2124_, new_n202_, new_n2165_})
4'b11?? : new_n2380_ = 1'b1;
4'b??10 : new_n2380_ = 1'b1;
default : new_n2380_ = 1'b0;
endcase
casez ({new_n1446_, new_n2226_})
2'b01 : new_n2381_ = 1'b1;
default : new_n2381_ = 1'b0;
endcase
casez ({new_n190_, new_n277_, new_n5921_})
3'b11? : new_n2382_ = 1'b1;
3'b??1 : new_n2382_ = 1'b1;
default : new_n2382_ = 1'b0;
endcase
casez ({new_n256_, new_n563_, new_n376_, new_n556_})
4'b11?? : new_n2383_ = 1'b1;
4'b??11 : new_n2383_ = 1'b1;
default : new_n2383_ = 1'b0;
endcase
casez ({new_n196_, new_n1290_, new_n445_, new_n562_})
4'b11?? : new_n2384_ = 1'b1;
4'b??11 : new_n2384_ = 1'b1;
default : new_n2384_ = 1'b0;
endcase
casez ({new_n144_, new_n415_, new_n346_, new_n876_})
4'b11?? : new_n2385_ = 1'b1;
4'b??11 : new_n2385_ = 1'b1;
default : new_n2385_ = 1'b0;
endcase
casez ({v[2], new_n879_, new_n268_, new_n618_})
4'b01?? : new_n2386_ = 1'b1;
4'b??11 : new_n2386_ = 1'b1;
default : new_n2386_ = 1'b0;
endcase
casez ({new_n88_, new_n585_, new_n5923_})
3'b11? : new_n2387_ = 1'b1;
3'b??1 : new_n2387_ = 1'b1;
default : new_n2387_ = 1'b0;
endcase
casez ({new_n728_, new_n3404_, new_n887_})
3'b11? : new_n2388_ = 1'b1;
3'b??1 : new_n2388_ = 1'b1;
default : new_n2388_ = 1'b0;
endcase
casez ({new_n129_, new_n685_, new_n139_, new_n892_})
4'b11?? : new_n2389_ = 1'b1;
4'b??11 : new_n2389_ = 1'b1;
default : new_n2389_ = 1'b0;
endcase
casez ({new_n304_, new_n894_, new_n597_, new_n802_})
4'b01?? : new_n2390_ = 1'b1;
4'b??11 : new_n2390_ = 1'b1;
default : new_n2390_ = 1'b0;
endcase
casez ({new_n182_, new_n560_, new_n355_, new_n1363_})
4'b11?? : new_n2391_ = 1'b1;
4'b??11 : new_n2391_ = 1'b1;
default : new_n2391_ = 1'b0;
endcase
casez ({new_n205_, new_n759_, new_n301_, new_n909_})
4'b10?? : new_n2392_ = 1'b1;
4'b??11 : new_n2392_ = 1'b1;
default : new_n2392_ = 1'b0;
endcase
casez ({new_n5924_, new_n305_, new_n915_})
3'b1?? : new_n2393_ = 1'b1;
3'b?11 : new_n2393_ = 1'b1;
default : new_n2393_ = 1'b0;
endcase
casez ({new_n691_, new_n1418_})
2'b00 : new_n2394_ = 1'b1;
default : new_n2394_ = 1'b0;
endcase
casez ({new_n664_, new_n1419_})
2'b00 : new_n2395_ = 1'b1;
default : new_n2395_ = 1'b0;
endcase
casez ({new_n174_, new_n589_, new_n194_, new_n1424_})
4'b11?? : new_n2396_ = 1'b1;
4'b??11 : new_n2396_ = 1'b1;
default : new_n2396_ = 1'b0;
endcase
casez ({new_n201_, new_n1439_, new_n310_, new_n1073_})
4'b11?? : new_n2397_ = 1'b1;
4'b??11 : new_n2397_ = 1'b1;
default : new_n2397_ = 1'b0;
endcase
casez ({new_n226_, new_n687_, new_n712_, new_n1440_})
4'b11?? : new_n2398_ = 1'b1;
4'b??11 : new_n2398_ = 1'b1;
default : new_n2398_ = 1'b0;
endcase
casez ({new_n792_, new_n1441_})
2'b00 : new_n2399_ = 1'b1;
default : new_n2399_ = 1'b0;
endcase
casez ({new_n182_, new_n1443_, new_n201_, new_n1106_})
4'b11?? : new_n2400_ = 1'b1;
4'b??11 : new_n2400_ = 1'b1;
default : new_n2400_ = 1'b0;
endcase
casez ({new_n88_, new_n1420_, new_n107_, new_n1451_})
4'b11?? : new_n2401_ = 1'b1;
4'b??01 : new_n2401_ = 1'b1;
default : new_n2401_ = 1'b0;
endcase
casez ({new_n885_, new_n1478_})
2'b00 : new_n2402_ = 1'b1;
default : new_n2402_ = 1'b0;
endcase
casez ({new_n588_, new_n1490_})
2'b00 : new_n2403_ = 1'b1;
default : new_n2403_ = 1'b0;
endcase
casez ({new_n255_, new_n1425_, new_n303_, new_n1514_})
4'b11?? : new_n2404_ = 1'b1;
4'b??10 : new_n2404_ = 1'b1;
default : new_n2404_ = 1'b0;
endcase
casez ({new_n161_, new_n640_, new_n171_, new_n1515_})
4'b11?? : new_n2405_ = 1'b1;
4'b??10 : new_n2405_ = 1'b1;
default : new_n2405_ = 1'b0;
endcase
casez ({new_n87_, new_n1526_, new_n456_, new_n501_})
4'b01?? : new_n2406_ = 1'b1;
4'b??11 : new_n2406_ = 1'b1;
default : new_n2406_ = 1'b0;
endcase
casez ({new_n158_, new_n547_, new_n366_, new_n653_})
4'b11?? : new_n2407_ = 1'b1;
4'b??11 : new_n2407_ = 1'b1;
default : new_n2407_ = 1'b0;
endcase
casez ({new_n916_, new_n1010_})
2'b00 : new_n2408_ = 1'b1;
default : new_n2408_ = 1'b0;
endcase
casez ({new_n390_, new_n990_, new_n429_, new_n1013_})
4'b11?? : new_n2409_ = 1'b1;
4'b??11 : new_n2409_ = 1'b1;
default : new_n2409_ = 1'b0;
endcase
casez ({new_n228_, new_n1021_, new_n377_, new_n622_})
4'b11?? : new_n2410_ = 1'b1;
4'b??11 : new_n2410_ = 1'b1;
default : new_n2410_ = 1'b0;
endcase
casez ({new_n155_, new_n688_, new_n240_, new_n569_})
4'b11?? : new_n2411_ = 1'b1;
4'b??11 : new_n2411_ = 1'b1;
default : new_n2411_ = 1'b0;
endcase
casez ({new_n122_, new_n690_, new_n164_, new_n587_})
4'b11?? : new_n2412_ = 1'b1;
4'b??11 : new_n2412_ = 1'b1;
default : new_n2412_ = 1'b0;
endcase
casez ({new_n176_, new_n643_, new_n221_, new_n1655_})
4'b11?? : new_n2413_ = 1'b1;
4'b??11 : new_n2413_ = 1'b1;
default : new_n2413_ = 1'b0;
endcase
casez ({new_n86_, new_n1459_, new_n150_, new_n1656_})
4'b11?? : new_n2414_ = 1'b1;
4'b??11 : new_n2414_ = 1'b1;
default : new_n2414_ = 1'b0;
endcase
casez ({new_n225_, new_n1657_, new_n607_, new_n727_})
4'b11?? : new_n2415_ = 1'b1;
4'b??11 : new_n2415_ = 1'b1;
default : new_n2415_ = 1'b0;
endcase
casez ({new_n1031_, new_n1658_})
2'b00 : new_n2416_ = 1'b1;
default : new_n2416_ = 1'b0;
endcase
casez ({new_n232_, new_n551_, new_n268_, new_n1052_})
4'b11?? : new_n2417_ = 1'b1;
4'b??11 : new_n2417_ = 1'b1;
default : new_n2417_ = 1'b0;
endcase
casez ({new_n139_, new_n1685_, new_n248_, new_n945_})
4'b11?? : new_n2418_ = 1'b1;
4'b??11 : new_n2418_ = 1'b1;
default : new_n2418_ = 1'b0;
endcase
casez ({new_n90_, new_n1695_, new_n91_, new_n1683_})
4'b11?? : new_n2419_ = 1'b1;
4'b??11 : new_n2419_ = 1'b1;
default : new_n2419_ = 1'b0;
endcase
casez ({new_n171_, new_n1698_, new_n347_, new_n810_})
4'b11?? : new_n2420_ = 1'b1;
4'b??11 : new_n2420_ = 1'b1;
default : new_n2420_ = 1'b0;
endcase
casez ({new_n340_, new_n1049_, new_n495_, new_n1707_})
4'b11?? : new_n2421_ = 1'b1;
4'b??11 : new_n2421_ = 1'b1;
default : new_n2421_ = 1'b0;
endcase
casez ({new_n155_, new_n890_, new_n250_, new_n1064_})
4'b11?? : new_n2422_ = 1'b1;
4'b??11 : new_n2422_ = 1'b1;
default : new_n2422_ = 1'b0;
endcase
casez ({new_n97_, new_n1614_, new_n148_, new_n1739_})
4'b11?? : new_n2423_ = 1'b1;
4'b??11 : new_n2423_ = 1'b1;
default : new_n2423_ = 1'b0;
endcase
casez ({new_n459_, new_n1073_, new_n916_, new_n927_})
4'b11?? : new_n2424_ = 1'b1;
4'b??11 : new_n2424_ = 1'b1;
default : new_n2424_ = 1'b0;
endcase
casez ({new_n396_, new_n452_})
2'b00 : new_n2425_ = 1'b1;
default : new_n2425_ = 1'b0;
endcase
casez ({new_n475_, new_n1114_})
2'b00 : new_n2426_ = 1'b1;
default : new_n2426_ = 1'b0;
endcase
casez ({new_n161_, new_n760_, new_n168_, new_n663_})
4'b11?? : new_n2427_ = 1'b1;
4'b??11 : new_n2427_ = 1'b1;
default : new_n2427_ = 1'b0;
endcase
casez ({new_n546_, new_n1819_, new_n1107_, new_n1888_})
4'b10?? : new_n2428_ = 1'b1;
4'b??11 : new_n2428_ = 1'b1;
default : new_n2428_ = 1'b0;
endcase
casez ({new_n117_, new_n169_})
2'b11 : new_n2429_ = 1'b1;
default : new_n2429_ = 1'b0;
endcase
casez ({new_n224_, new_n1085_, new_n906_, new_n1161_})
4'b11?? : new_n2430_ = 1'b1;
4'b??11 : new_n2430_ = 1'b1;
default : new_n2430_ = 1'b0;
endcase
casez ({new_n187_, new_n374_, new_n416_, new_n793_})
4'b11?? : new_n2431_ = 1'b1;
4'b??11 : new_n2431_ = 1'b1;
default : new_n2431_ = 1'b0;
endcase
casez ({new_n331_, new_n2974_, new_n2009_})
3'b11? : new_n2432_ = 1'b1;
3'b??1 : new_n2432_ = 1'b1;
default : new_n2432_ = 1'b0;
endcase
casez ({new_n353_, new_n3451_, new_n1230_})
3'b11? : new_n2433_ = 1'b1;
3'b??1 : new_n2433_ = 1'b1;
default : new_n2433_ = 1'b0;
endcase
casez ({new_n212_, new_n4615_, new_n1231_})
3'b11? : new_n2434_ = 1'b1;
3'b??1 : new_n2434_ = 1'b1;
default : new_n2434_ = 1'b0;
endcase
casez ({v[0], new_n273_, new_n680_, new_n1235_})
4'b111? : new_n2435_ = 1'b1;
4'b???1 : new_n2435_ = 1'b1;
default : new_n2435_ = 1'b0;
endcase
casez ({new_n253_, new_n3464_, new_n2169_})
3'b11? : new_n2436_ = 1'b1;
3'b??1 : new_n2436_ = 1'b1;
default : new_n2436_ = 1'b0;
endcase
casez ({new_n87_, new_n120_, new_n542_, new_n2178_})
4'b111? : new_n2437_ = 1'b1;
4'b???1 : new_n2437_ = 1'b1;
default : new_n2437_ = 1'b0;
endcase
casez ({new_n4618_, new_n2180_})
2'b1? : new_n2438_ = 1'b1;
2'b?1 : new_n2438_ = 1'b1;
default : new_n2438_ = 1'b0;
endcase
casez ({new_n184_, new_n226_, new_n249_, new_n2181_})
4'b111? : new_n2439_ = 1'b1;
4'b???1 : new_n2439_ = 1'b1;
default : new_n2439_ = 1'b0;
endcase
casez ({new_n104_, new_n207_, new_n606_, new_n2203_})
4'b111? : new_n2440_ = 1'b1;
4'b???1 : new_n2440_ = 1'b1;
default : new_n2440_ = 1'b0;
endcase
casez ({new_n346_, new_n3531_, new_n2206_})
3'b11? : new_n2441_ = 1'b1;
3'b??1 : new_n2441_ = 1'b1;
default : new_n2441_ = 1'b0;
endcase
casez ({new_n786_, new_n3576_, new_n2208_})
3'b11? : new_n2442_ = 1'b1;
3'b??1 : new_n2442_ = 1'b1;
default : new_n2442_ = 1'b0;
endcase
casez ({new_n226_, new_n3395_, new_n2216_})
3'b11? : new_n2443_ = 1'b1;
3'b??1 : new_n2443_ = 1'b1;
default : new_n2443_ = 1'b0;
endcase
casez ({v[0], new_n97_, new_n1265_, new_n1239_})
4'b011? : new_n2444_ = 1'b1;
4'b???1 : new_n2444_ = 1'b1;
default : new_n2444_ = 1'b0;
endcase
casez ({new_n338_, new_n4619_, new_n2220_})
3'b11? : new_n2445_ = 1'b1;
3'b??1 : new_n2445_ = 1'b1;
default : new_n2445_ = 1'b0;
endcase
casez ({y[2], new_n100_, new_n1744_, new_n2223_})
4'b011? : new_n2446_ = 1'b1;
4'b???1 : new_n2446_ = 1'b1;
default : new_n2446_ = 1'b0;
endcase
casez ({new_n495_, new_n3573_, new_n2229_})
3'b11? : new_n2447_ = 1'b1;
3'b??1 : new_n2447_ = 1'b1;
default : new_n2447_ = 1'b0;
endcase
casez ({new_n623_, new_n3472_, new_n2231_})
3'b11? : new_n2448_ = 1'b1;
3'b??1 : new_n2448_ = 1'b1;
default : new_n2448_ = 1'b0;
endcase
casez ({new_n84_, new_n386_, new_n414_, new_n2257_})
4'b111? : new_n2449_ = 1'b1;
4'b???1 : new_n2449_ = 1'b1;
default : new_n2449_ = 1'b0;
endcase
casez ({new_n906_, new_n3346_, new_n2263_})
3'b11? : new_n2450_ = 1'b1;
3'b??1 : new_n2450_ = 1'b1;
default : new_n2450_ = 1'b0;
endcase
casez ({v[1], new_n240_, new_n334_, new_n2264_})
4'b011? : new_n2451_ = 1'b1;
4'b???1 : new_n2451_ = 1'b1;
default : new_n2451_ = 1'b0;
endcase
casez ({new_n112_, new_n3457_, new_n2278_})
3'b11? : new_n2452_ = 1'b1;
3'b??1 : new_n2452_ = 1'b1;
default : new_n2452_ = 1'b0;
endcase
casez ({new_n132_, new_n150_, new_n258_, new_n2290_})
4'b111? : new_n2453_ = 1'b1;
4'b???1 : new_n2453_ = 1'b1;
default : new_n2453_ = 1'b0;
endcase
casez ({new_n140_, new_n278_, new_n287_, new_n2294_})
4'b111? : new_n2454_ = 1'b1;
4'b???1 : new_n2454_ = 1'b1;
default : new_n2454_ = 1'b0;
endcase
casez ({new_n154_, new_n3354_, new_n2305_})
3'b11? : new_n2455_ = 1'b1;
3'b??1 : new_n2455_ = 1'b1;
default : new_n2455_ = 1'b0;
endcase
casez ({new_n508_, new_n3551_, new_n2308_})
3'b11? : new_n2456_ = 1'b1;
3'b??1 : new_n2456_ = 1'b1;
default : new_n2456_ = 1'b0;
endcase
casez ({new_n120_, new_n4622_, new_n2319_})
3'b11? : new_n2457_ = 1'b1;
3'b??1 : new_n2457_ = 1'b1;
default : new_n2457_ = 1'b0;
endcase
casez ({new_n304_, new_n1079_, new_n406_, new_n2381_})
4'b01?? : new_n2458_ = 1'b1;
4'b??00 : new_n2458_ = 1'b1;
default : new_n2458_ = 1'b0;
endcase
casez ({new_n160_, new_n2394_, new_n219_, new_n1677_})
4'b10?? : new_n2459_ = 1'b1;
4'b??11 : new_n2459_ = 1'b1;
default : new_n2459_ = 1'b0;
endcase
casez ({new_n113_, new_n1084_, new_n298_, new_n1398_})
4'b11?? : new_n2460_ = 1'b1;
4'b??11 : new_n2460_ = 1'b1;
default : new_n2460_ = 1'b0;
endcase
casez ({new_n81_, new_n1432_, new_n6128_})
3'b11? : new_n2461_ = 1'b1;
3'b??1 : new_n2461_ = 1'b1;
default : new_n2461_ = 1'b0;
endcase
casez ({new_n167_, new_n700_, new_n478_, new_n1467_})
4'b11?? : new_n2462_ = 1'b1;
4'b??11 : new_n2462_ = 1'b1;
default : new_n2462_ = 1'b0;
endcase
casez ({new_n183_, new_n375_, new_n213_, new_n1512_})
4'b11?? : new_n2463_ = 1'b1;
4'b??11 : new_n2463_ = 1'b1;
default : new_n2463_ = 1'b0;
endcase
casez ({new_n90_, new_n1523_, new_n375_, new_n709_})
4'b11?? : new_n2464_ = 1'b1;
4'b??10 : new_n2464_ = 1'b1;
default : new_n2464_ = 1'b0;
endcase
casez ({new_n168_, new_n1534_, new_n176_, new_n1004_})
4'b10?? : new_n2465_ = 1'b1;
4'b??11 : new_n2465_ = 1'b1;
default : new_n2465_ = 1'b0;
endcase
casez ({new_n396_, new_n1535_, new_n441_, new_n1521_})
4'b10?? : new_n2466_ = 1'b1;
4'b??11 : new_n2466_ = 1'b1;
default : new_n2466_ = 1'b0;
endcase
casez ({new_n214_, new_n1036_, new_n262_, new_n762_})
4'b11?? : new_n2467_ = 1'b1;
4'b??11 : new_n2467_ = 1'b1;
default : new_n2467_ = 1'b0;
endcase
casez ({new_n149_, new_n327_, new_n375_, new_n403_})
4'b11?? : new_n2468_ = 1'b1;
4'b??11 : new_n2468_ = 1'b1;
default : new_n2468_ = 1'b0;
endcase
casez ({new_n211_, new_n1518_, new_n554_, new_n1662_})
4'b11?? : new_n2469_ = 1'b1;
4'b??11 : new_n2469_ = 1'b1;
default : new_n2469_ = 1'b0;
endcase
casez ({new_n82_, new_n762_, new_n183_, new_n1078_})
4'b11?? : new_n2470_ = 1'b1;
4'b??11 : new_n2470_ = 1'b1;
default : new_n2470_ = 1'b0;
endcase
casez ({new_n89_, new_n1511_, new_n288_, new_n1767_})
4'b11?? : new_n2471_ = 1'b1;
4'b??01 : new_n2471_ = 1'b1;
default : new_n2471_ = 1'b0;
endcase
casez ({new_n101_, new_n294_, new_n332_, new_n1788_})
4'b111? : new_n2472_ = 1'b1;
4'b???1 : new_n2472_ = 1'b1;
default : new_n2472_ = 1'b0;
endcase
casez ({new_n594_, new_n738_})
2'b00 : new_n2473_ = 1'b1;
default : new_n2473_ = 1'b0;
endcase
casez ({new_n305_, new_n626_, new_n375_, new_n752_})
4'b11?? : new_n2474_ = 1'b1;
4'b??11 : new_n2474_ = 1'b1;
default : new_n2474_ = 1'b0;
endcase
casez ({new_n116_, new_n375_, new_n171_, new_n474_})
4'b11?? : new_n2475_ = 1'b1;
4'b??11 : new_n2475_ = 1'b1;
default : new_n2475_ = 1'b0;
endcase
casez ({new_n95_, new_n96_, new_n950_, new_n1248_})
4'b111? : new_n2476_ = 1'b1;
4'b???1 : new_n2476_ = 1'b1;
default : new_n2476_ = 1'b0;
endcase
casez ({new_n672_, new_n3483_, new_n2358_})
3'b11? : new_n2477_ = 1'b1;
3'b??1 : new_n2477_ = 1'b1;
default : new_n2477_ = 1'b0;
endcase
casez ({new_n4608_, new_n2370_})
2'b1? : new_n2478_ = 1'b1;
2'b?1 : new_n2478_ = 1'b1;
default : new_n2478_ = 1'b0;
endcase
casez ({new_n355_, new_n3492_, new_n2380_})
3'b11? : new_n2479_ = 1'b1;
3'b??1 : new_n2479_ = 1'b1;
default : new_n2479_ = 1'b0;
endcase
casez ({new_n98_, new_n100_, new_n730_, new_n2382_})
4'b111? : new_n2480_ = 1'b1;
4'b???1 : new_n2480_ = 1'b1;
default : new_n2480_ = 1'b0;
endcase
casez ({new_n142_, new_n4593_, new_n2384_})
3'b11? : new_n2481_ = 1'b1;
3'b??1 : new_n2481_ = 1'b1;
default : new_n2481_ = 1'b0;
endcase
casez ({new_n118_, new_n127_, new_n200_, new_n2418_})
4'b111? : new_n2482_ = 1'b1;
4'b???1 : new_n2482_ = 1'b1;
default : new_n2482_ = 1'b0;
endcase
casez ({new_n218_, new_n820_, new_n1002_, new_n1397_})
4'b11?? : new_n2483_ = 1'b1;
4'b??11 : new_n2483_ = 1'b1;
default : new_n2483_ = 1'b0;
endcase
casez ({new_n228_, new_n614_, new_n286_, new_n375_})
4'b11?? : new_n2484_ = 1'b1;
4'b??11 : new_n2484_ = 1'b1;
default : new_n2484_ = 1'b0;
endcase
casez ({u[0], new_n456_, new_n1189_, new_n1527_})
4'b011? : new_n2485_ = 1'b1;
4'b???1 : new_n2485_ = 1'b1;
default : new_n2485_ = 1'b0;
endcase
casez ({new_n84_, new_n1532_, new_n431_, new_n1531_})
4'b11?? : new_n2486_ = 1'b1;
4'b??11 : new_n2486_ = 1'b1;
default : new_n2486_ = 1'b0;
endcase
casez ({new_n158_, new_n1081_, new_n171_, new_n820_})
4'b11?? : new_n2487_ = 1'b1;
4'b??11 : new_n2487_ = 1'b1;
default : new_n2487_ = 1'b0;
endcase
casez ({new_n217_, new_n1089_, new_n375_, new_n454_})
4'b11?? : new_n2488_ = 1'b1;
4'b??11 : new_n2488_ = 1'b1;
default : new_n2488_ = 1'b0;
endcase
casez ({new_n266_, new_n1089_, new_n499_, new_n614_})
4'b11?? : new_n2489_ = 1'b1;
4'b??11 : new_n2489_ = 1'b1;
default : new_n2489_ = 1'b0;
endcase
casez ({new_n82_, new_n1784_, new_n5925_})
3'b11? : new_n2490_ = 1'b1;
3'b??1 : new_n2490_ = 1'b1;
default : new_n2490_ = 1'b0;
endcase
casez ({new_n363_, new_n3410_, new_n2430_})
3'b11? : new_n2491_ = 1'b1;
3'b??1 : new_n2491_ = 1'b1;
default : new_n2491_ = 1'b0;
endcase
casez ({new_n400_, new_n1756_, new_n574_, new_n1538_})
4'b11?? : new_n2492_ = 1'b1;
4'b??01 : new_n2492_ = 1'b1;
default : new_n2492_ = 1'b0;
endcase
casez ({new_n260_, new_n1774_, new_n507_, new_n2379_})
4'b11?? : new_n2493_ = 1'b1;
4'b??10 : new_n2493_ = 1'b1;
default : new_n2493_ = 1'b0;
endcase
casez ({new_n456_, new_n3456_, new_n922_})
3'b11? : new_n2494_ = 1'b1;
3'b??1 : new_n2494_ = 1'b1;
default : new_n2494_ = 1'b0;
endcase
casez ({y[1], v[0]})
2'b10 : new_n2495_ = 1'b1;
default : new_n2495_ = 1'b0;
endcase
casez ({x[2], u[2]})
2'b11 : new_n2496_ = 1'b1;
default : new_n2496_ = 1'b0;
endcase
casez ({x[0], u[1]})
2'b11 : new_n2497_ = 1'b1;
default : new_n2497_ = 1'b0;
endcase
casez ({x[1], v[1], new_n98_})
3'b00? : new_n2498_ = 1'b1;
3'b??1 : new_n2498_ = 1'b1;
default : new_n2498_ = 1'b0;
endcase
casez ({new_n2939_, new_n98_})
2'b1? : new_n2499_ = 1'b1;
2'b?1 : new_n2499_ = 1'b1;
default : new_n2499_ = 1'b0;
endcase
casez ({new_n84_, new_n328_})
2'b00 : new_n2500_ = 1'b1;
default : new_n2500_ = 1'b0;
endcase
casez ({v[1], new_n92_})
2'b11 : new_n2501_ = 1'b1;
default : new_n2501_ = 1'b0;
endcase
casez ({u[2], new_n104_})
2'b01 : new_n2502_ = 1'b1;
default : new_n2502_ = 1'b0;
endcase
casez ({new_n86_, new_n89_})
2'b10 : new_n2503_ = 1'b1;
default : new_n2503_ = 1'b0;
endcase
casez ({new_n82_, new_n90_})
2'b10 : new_n2504_ = 1'b1;
default : new_n2504_ = 1'b0;
endcase
casez ({new_n81_, new_n90_})
2'b10 : new_n2505_ = 1'b1;
default : new_n2505_ = 1'b0;
endcase
casez ({x[1], new_n278_})
2'b11 : new_n2506_ = 1'b1;
default : new_n2506_ = 1'b0;
endcase
casez ({new_n80_, new_n281_})
2'b11 : new_n2507_ = 1'b1;
default : new_n2507_ = 1'b0;
endcase
casez ({x[1], new_n281_})
2'b01 : new_n2508_ = 1'b1;
default : new_n2508_ = 1'b0;
endcase
casez ({y[0], new_n94_})
2'b00 : new_n2509_ = 1'b1;
default : new_n2509_ = 1'b0;
endcase
casez ({new_n90_, new_n94_})
2'b01 : new_n2510_ = 1'b1;
default : new_n2510_ = 1'b0;
endcase
casez ({new_n91_, new_n95_})
2'b01 : new_n2511_ = 1'b1;
default : new_n2511_ = 1'b0;
endcase
casez ({new_n97_, new_n315_})
2'b11 : new_n2512_ = 1'b1;
default : new_n2512_ = 1'b0;
endcase
casez ({new_n82_, new_n100_})
2'b10 : new_n2513_ = 1'b1;
default : new_n2513_ = 1'b0;
endcase
casez ({v[2], new_n100_})
2'b00 : new_n2514_ = 1'b1;
default : new_n2514_ = 1'b0;
endcase
casez ({new_n88_, new_n104_})
2'b10 : new_n2515_ = 1'b1;
default : new_n2515_ = 1'b0;
endcase
casez ({new_n80_, new_n385_})
2'b11 : new_n2516_ = 1'b1;
default : new_n2516_ = 1'b0;
endcase
casez ({new_n91_, new_n94_})
2'b01 : new_n2517_ = 1'b1;
default : new_n2517_ = 1'b0;
endcase
casez ({new_n94_, new_n100_})
2'b10 : new_n2518_ = 1'b1;
default : new_n2518_ = 1'b0;
endcase
casez ({new_n80_, new_n88_})
2'b11 : new_n2519_ = 1'b1;
default : new_n2519_ = 1'b0;
endcase
casez ({new_n89_, new_n93_})
2'b11 : new_n2520_ = 1'b1;
default : new_n2520_ = 1'b0;
endcase
casez ({new_n86_, new_n93_})
2'b11 : new_n2521_ = 1'b1;
default : new_n2521_ = 1'b0;
endcase
casez ({y[0], new_n98_})
2'b11 : new_n2522_ = 1'b1;
default : new_n2522_ = 1'b0;
endcase
casez ({new_n191_, new_n251_})
2'b00 : new_n2523_ = 1'b1;
default : new_n2523_ = 1'b0;
endcase
casez ({new_n95_, new_n100_, new_n255_})
3'b10? : new_n2524_ = 1'b1;
3'b??1 : new_n2524_ = 1'b1;
default : new_n2524_ = 1'b0;
endcase
casez ({new_n115_, new_n150_})
2'b00 : new_n2525_ = 1'b1;
default : new_n2525_ = 1'b0;
endcase
casez ({new_n161_, new_n278_})
2'b00 : new_n2526_ = 1'b1;
default : new_n2526_ = 1'b0;
endcase
casez ({new_n103_, new_n159_})
2'b00 : new_n2527_ = 1'b1;
default : new_n2527_ = 1'b0;
endcase
casez ({new_n158_, new_n160_})
2'b00 : new_n2528_ = 1'b1;
default : new_n2528_ = 1'b0;
endcase
casez ({new_n116_, new_n163_})
2'b00 : new_n2529_ = 1'b1;
default : new_n2529_ = 1'b0;
endcase
casez ({new_n204_, new_n1261_})
2'b01 : new_n2530_ = 1'b1;
default : new_n2530_ = 1'b0;
endcase
casez ({new_n210_, new_n301_})
2'b00 : new_n2531_ = 1'b1;
default : new_n2531_ = 1'b0;
endcase
casez ({new_n159_, new_n177_})
2'b00 : new_n2532_ = 1'b1;
default : new_n2532_ = 1'b0;
endcase
casez ({new_n211_, new_n317_})
2'b00 : new_n2533_ = 1'b1;
default : new_n2533_ = 1'b0;
endcase
casez ({new_n235_, new_n2517_})
2'b00 : new_n2534_ = 1'b1;
default : new_n2534_ = 1'b0;
endcase
casez ({new_n198_, new_n321_})
2'b00 : new_n2535_ = 1'b1;
default : new_n2535_ = 1'b0;
endcase
casez ({new_n183_, new_n184_})
2'b00 : new_n2536_ = 1'b1;
default : new_n2536_ = 1'b0;
endcase
casez ({new_n239_, new_n927_})
2'b00 : new_n2537_ = 1'b1;
default : new_n2537_ = 1'b0;
endcase
casez ({new_n213_, new_n342_})
2'b00 : new_n2538_ = 1'b1;
default : new_n2538_ = 1'b0;
endcase
casez ({new_n293_, new_n344_})
2'b00 : new_n2539_ = 1'b1;
default : new_n2539_ = 1'b0;
endcase
casez ({new_n293_, new_n347_})
2'b00 : new_n2540_ = 1'b1;
default : new_n2540_ = 1'b0;
endcase
casez ({new_n167_, new_n347_})
2'b00 : new_n2541_ = 1'b1;
default : new_n2541_ = 1'b0;
endcase
casez ({new_n159_, new_n199_})
2'b00 : new_n2542_ = 1'b1;
default : new_n2542_ = 1'b0;
endcase
casez ({new_n192_, new_n199_})
2'b00 : new_n2543_ = 1'b1;
default : new_n2543_ = 1'b0;
endcase
casez ({new_n158_, new_n201_})
2'b00 : new_n2544_ = 1'b1;
default : new_n2544_ = 1'b0;
endcase
casez ({new_n178_, new_n208_})
2'b00 : new_n2545_ = 1'b1;
default : new_n2545_ = 1'b0;
endcase
casez ({new_n192_, new_n208_})
2'b00 : new_n2546_ = 1'b1;
default : new_n2546_ = 1'b0;
endcase
casez ({new_n167_, new_n215_})
2'b00 : new_n2547_ = 1'b1;
default : new_n2547_ = 1'b0;
endcase
casez ({new_n155_, new_n218_})
2'b00 : new_n2548_ = 1'b1;
default : new_n2548_ = 1'b0;
endcase
casez ({new_n190_, new_n226_})
2'b00 : new_n2549_ = 1'b1;
default : new_n2549_ = 1'b0;
endcase
casez ({new_n90_, new_n228_})
2'b00 : new_n2550_ = 1'b1;
default : new_n2550_ = 1'b0;
endcase
casez ({new_n77_, new_n437_})
2'b00 : new_n2551_ = 1'b1;
default : new_n2551_ = 1'b0;
endcase
casez ({new_n221_, new_n240_})
2'b00 : new_n2552_ = 1'b1;
default : new_n2552_ = 1'b0;
endcase
casez ({v[0], new_n77_})
2'b11 : new_n2553_ = 1'b1;
default : new_n2553_ = 1'b0;
endcase
casez ({new_n243_, new_n254_})
2'b11 : new_n2554_ = 1'b1;
default : new_n2554_ = 1'b0;
endcase
casez ({new_n162_, new_n255_})
2'b11 : new_n2555_ = 1'b1;
default : new_n2555_ = 1'b0;
endcase
casez ({new_n234_, new_n488_})
2'b11 : new_n2556_ = 1'b1;
default : new_n2556_ = 1'b0;
endcase
casez ({new_n207_, new_n255_})
2'b11 : new_n2557_ = 1'b1;
default : new_n2557_ = 1'b0;
endcase
casez ({new_n144_, new_n488_})
2'b11 : new_n2558_ = 1'b1;
default : new_n2558_ = 1'b0;
endcase
casez ({new_n344_, new_n489_})
2'b11 : new_n2559_ = 1'b1;
default : new_n2559_ = 1'b0;
endcase
casez ({new_n118_, new_n254_})
2'b11 : new_n2560_ = 1'b1;
default : new_n2560_ = 1'b0;
endcase
casez ({new_n137_, new_n258_})
2'b11 : new_n2561_ = 1'b1;
default : new_n2561_ = 1'b0;
endcase
casez ({new_n209_, new_n258_})
2'b11 : new_n2562_ = 1'b1;
default : new_n2562_ = 1'b0;
endcase
casez ({new_n167_, new_n262_})
2'b11 : new_n2563_ = 1'b1;
default : new_n2563_ = 1'b0;
endcase
casez ({new_n248_, new_n262_})
2'b11 : new_n2564_ = 1'b1;
default : new_n2564_ = 1'b0;
endcase
casez ({new_n234_, new_n508_})
2'b11 : new_n2565_ = 1'b1;
default : new_n2565_ = 1'b0;
endcase
casez ({new_n228_, new_n2565_, new_n1599_, new_n2495_})
4'b11?? : new_n2566_ = 1'b1;
4'b??11 : new_n2566_ = 1'b1;
default : new_n2566_ = 1'b0;
endcase
casez ({x[1], new_n1090_, new_n1613_, new_n2566_})
4'b011? : new_n2567_ = 1'b1;
4'b???1 : new_n2567_ = 1'b1;
default : new_n2567_ = 1'b0;
endcase
casez ({new_n145_, new_n148_})
2'b11 : new_n2568_ = 1'b1;
default : new_n2568_ = 1'b0;
endcase
casez ({new_n176_, new_n273_})
2'b11 : new_n2569_ = 1'b1;
default : new_n2569_ = 1'b0;
endcase
casez ({new_n173_, new_n2569_, new_n290_, new_n1848_})
4'b11?? : new_n2570_ = 1'b1;
4'b??11 : new_n2570_ = 1'b1;
default : new_n2570_ = 1'b0;
endcase
casez ({new_n155_, new_n273_})
2'b11 : new_n2571_ = 1'b1;
default : new_n2571_ = 1'b0;
endcase
casez ({new_n166_, new_n275_})
2'b11 : new_n2572_ = 1'b1;
default : new_n2572_ = 1'b0;
endcase
casez ({new_n224_, new_n275_})
2'b11 : new_n2573_ = 1'b1;
default : new_n2573_ = 1'b0;
endcase
casez ({new_n145_, new_n158_})
2'b11 : new_n2574_ = 1'b1;
default : new_n2574_ = 1'b0;
endcase
casez ({new_n118_, new_n279_})
2'b11 : new_n2575_ = 1'b1;
default : new_n2575_ = 1'b0;
endcase
casez ({new_n131_, new_n160_})
2'b11 : new_n2576_ = 1'b1;
default : new_n2576_ = 1'b0;
endcase
casez ({new_n151_, new_n162_})
2'b11 : new_n2577_ = 1'b1;
default : new_n2577_ = 1'b0;
endcase
casez ({new_n159_, new_n162_})
2'b11 : new_n2578_ = 1'b1;
default : new_n2578_ = 1'b0;
endcase
casez ({new_n150_, new_n284_})
2'b11 : new_n2579_ = 1'b1;
default : new_n2579_ = 1'b0;
endcase
casez ({new_n139_, new_n284_})
2'b11 : new_n2580_ = 1'b1;
default : new_n2580_ = 1'b0;
endcase
casez ({new_n207_, new_n285_})
2'b11 : new_n2581_ = 1'b1;
default : new_n2581_ = 1'b0;
endcase
casez ({new_n77_, new_n165_})
2'b01 : new_n2582_ = 1'b1;
default : new_n2582_ = 1'b0;
endcase
casez ({y[1], new_n165_})
2'b01 : new_n2583_ = 1'b1;
default : new_n2583_ = 1'b0;
endcase
casez ({x[2], new_n287_})
2'b01 : new_n2584_ = 1'b1;
default : new_n2584_ = 1'b0;
endcase
casez ({new_n215_, new_n287_})
2'b11 : new_n2585_ = 1'b1;
default : new_n2585_ = 1'b0;
endcase
casez ({new_n616_, new_n1265_})
2'b11 : new_n2586_ = 1'b1;
default : new_n2586_ = 1'b0;
endcase
casez ({new_n129_, new_n169_})
2'b11 : new_n2587_ = 1'b1;
default : new_n2587_ = 1'b0;
endcase
casez ({new_n215_, new_n299_})
2'b11 : new_n2588_ = 1'b1;
default : new_n2588_ = 1'b0;
endcase
casez ({new_n191_, new_n274_})
2'b11 : new_n2589_ = 1'b1;
default : new_n2589_ = 1'b0;
endcase
casez ({new_n150_, new_n151_})
2'b11 : new_n2590_ = 1'b1;
default : new_n2590_ = 1'b0;
endcase
casez ({new_n139_, new_n176_})
2'b11 : new_n2591_ = 1'b1;
default : new_n2591_ = 1'b0;
endcase
casez ({new_n79_, new_n176_})
2'b01 : new_n2592_ = 1'b1;
default : new_n2592_ = 1'b0;
endcase
casez ({new_n85_, new_n309_})
2'b11 : new_n2593_ = 1'b1;
default : new_n2593_ = 1'b0;
endcase
casez ({new_n104_, new_n309_})
2'b11 : new_n2594_ = 1'b1;
default : new_n2594_ = 1'b0;
endcase
casez ({new_n151_, new_n309_})
2'b11 : new_n2595_ = 1'b1;
default : new_n2595_ = 1'b0;
endcase
casez ({new_n142_, new_n177_})
2'b11 : new_n2596_ = 1'b1;
default : new_n2596_ = 1'b0;
endcase
casez ({new_n144_, new_n509_})
2'b11 : new_n2597_ = 1'b1;
default : new_n2597_ = 1'b0;
endcase
casez ({new_n196_, new_n316_})
2'b11 : new_n2598_ = 1'b1;
default : new_n2598_ = 1'b0;
endcase
casez ({v[2], new_n180_})
2'b01 : new_n2599_ = 1'b1;
default : new_n2599_ = 1'b0;
endcase
casez ({new_n115_, new_n301_})
2'b11 : new_n2600_ = 1'b1;
default : new_n2600_ = 1'b0;
endcase
casez ({new_n209_, new_n301_})
2'b11 : new_n2601_ = 1'b1;
default : new_n2601_ = 1'b0;
endcase
casez ({new_n167_, new_n316_})
2'b11 : new_n2602_ = 1'b1;
default : new_n2602_ = 1'b0;
endcase
casez ({new_n123_, new_n321_})
2'b11 : new_n2603_ = 1'b1;
default : new_n2603_ = 1'b0;
endcase
casez ({new_n189_, new_n321_})
2'b11 : new_n2604_ = 1'b1;
default : new_n2604_ = 1'b0;
endcase
casez ({new_n137_, new_n328_})
2'b11 : new_n2605_ = 1'b1;
default : new_n2605_ = 1'b0;
endcase
casez ({new_n173_, new_n328_})
2'b11 : new_n2606_ = 1'b1;
default : new_n2606_ = 1'b0;
endcase
casez ({new_n150_, new_n926_})
2'b11 : new_n2607_ = 1'b1;
default : new_n2607_ = 1'b0;
endcase
casez ({new_n145_, new_n305_})
2'b11 : new_n2608_ = 1'b1;
default : new_n2608_ = 1'b0;
endcase
casez ({new_n155_, new_n332_})
2'b11 : new_n2609_ = 1'b1;
default : new_n2609_ = 1'b0;
endcase
casez ({new_n162_, new_n189_})
2'b11 : new_n2610_ = 1'b1;
default : new_n2610_ = 1'b0;
endcase
casez ({new_n97_, new_n190_})
2'b01 : new_n2611_ = 1'b1;
default : new_n2611_ = 1'b0;
endcase
casez ({new_n142_, new_n190_})
2'b11 : new_n2612_ = 1'b1;
default : new_n2612_ = 1'b0;
endcase
casez ({new_n151_, new_n338_})
2'b11 : new_n2613_ = 1'b1;
default : new_n2613_ = 1'b0;
endcase
casez ({new_n166_, new_n338_})
2'b11 : new_n2614_ = 1'b1;
default : new_n2614_ = 1'b0;
endcase
casez ({new_n191_, new_n194_})
2'b11 : new_n2615_ = 1'b1;
default : new_n2615_ = 1'b0;
endcase
casez ({new_n170_, new_n194_})
2'b11 : new_n2616_ = 1'b1;
default : new_n2616_ = 1'b0;
endcase
casez ({u[1], new_n343_})
2'b01 : new_n2617_ = 1'b1;
default : new_n2617_ = 1'b0;
endcase
casez ({new_n224_, new_n343_})
2'b11 : new_n2618_ = 1'b1;
default : new_n2618_ = 1'b0;
endcase
casez ({new_n242_, new_n343_})
2'b11 : new_n2619_ = 1'b1;
default : new_n2619_ = 1'b0;
endcase
casez ({new_n107_, new_n196_})
2'b01 : new_n2620_ = 1'b1;
default : new_n2620_ = 1'b0;
endcase
casez ({new_n93_, new_n344_})
2'b11 : new_n2621_ = 1'b1;
default : new_n2621_ = 1'b0;
endcase
casez ({new_n182_, new_n198_})
2'b11 : new_n2622_ = 1'b1;
default : new_n2622_ = 1'b0;
endcase
casez ({new_n150_, new_n200_})
2'b11 : new_n2623_ = 1'b1;
default : new_n2623_ = 1'b0;
endcase
casez ({new_n248_, new_n351_})
2'b11 : new_n2624_ = 1'b1;
default : new_n2624_ = 1'b0;
endcase
casez ({new_n97_, new_n351_})
2'b11 : new_n2625_ = 1'b1;
default : new_n2625_ = 1'b0;
endcase
casez ({new_n177_, new_n356_})
2'b11 : new_n2626_ = 1'b1;
default : new_n2626_ = 1'b0;
endcase
casez ({new_n160_, new_n356_})
2'b11 : new_n2627_ = 1'b1;
default : new_n2627_ = 1'b0;
endcase
casez ({new_n176_, new_n358_})
2'b11 : new_n2628_ = 1'b1;
default : new_n2628_ = 1'b0;
endcase
casez ({new_n254_, new_n358_})
2'b11 : new_n2629_ = 1'b1;
default : new_n2629_ = 1'b0;
endcase
casez ({v[1], new_n205_})
2'b01 : new_n2630_ = 1'b1;
default : new_n2630_ = 1'b0;
endcase
casez ({new_n166_, new_n363_})
2'b11 : new_n2631_ = 1'b1;
default : new_n2631_ = 1'b0;
endcase
casez ({y[0], new_n654_})
2'b11 : new_n2632_ = 1'b1;
default : new_n2632_ = 1'b0;
endcase
casez ({new_n150_, new_n208_})
2'b11 : new_n2633_ = 1'b1;
default : new_n2633_ = 1'b0;
endcase
casez ({new_n201_, new_n369_})
2'b11 : new_n2634_ = 1'b1;
default : new_n2634_ = 1'b0;
endcase
casez ({new_n92_, new_n208_})
2'b01 : new_n2635_ = 1'b1;
default : new_n2635_ = 1'b0;
endcase
casez ({new_n167_, new_n209_})
2'b11 : new_n2636_ = 1'b1;
default : new_n2636_ = 1'b0;
endcase
casez ({new_n176_, new_n209_})
2'b11 : new_n2637_ = 1'b1;
default : new_n2637_ = 1'b0;
endcase
casez ({new_n118_, new_n210_})
2'b11 : new_n2638_ = 1'b1;
default : new_n2638_ = 1'b0;
endcase
casez ({new_n86_, new_n211_})
2'b01 : new_n2639_ = 1'b1;
default : new_n2639_ = 1'b0;
endcase
casez ({new_n166_, new_n211_})
2'b11 : new_n2640_ = 1'b1;
default : new_n2640_ = 1'b0;
endcase
casez ({new_n191_, new_n211_})
2'b11 : new_n2641_ = 1'b1;
default : new_n2641_ = 1'b0;
endcase
casez ({new_n184_, new_n212_})
2'b11 : new_n2642_ = 1'b1;
default : new_n2642_ = 1'b0;
endcase
casez ({new_n176_, new_n212_})
2'b11 : new_n2643_ = 1'b1;
default : new_n2643_ = 1'b0;
endcase
casez ({new_n150_, new_n385_})
2'b11 : new_n2644_ = 1'b1;
default : new_n2644_ = 1'b0;
endcase
casez ({new_n170_, new_n214_})
2'b11 : new_n2645_ = 1'b1;
default : new_n2645_ = 1'b0;
endcase
casez ({new_n189_, new_n216_})
2'b11 : new_n2646_ = 1'b1;
default : new_n2646_ = 1'b0;
endcase
casez ({new_n161_, new_n216_})
2'b11 : new_n2647_ = 1'b1;
default : new_n2647_ = 1'b0;
endcase
casez ({new_n215_, new_n219_})
2'b11 : new_n2648_ = 1'b1;
default : new_n2648_ = 1'b0;
endcase
casez ({new_n160_, new_n219_})
2'b11 : new_n2649_ = 1'b1;
default : new_n2649_ = 1'b0;
endcase
casez ({new_n170_, new_n219_})
2'b11 : new_n2650_ = 1'b1;
default : new_n2650_ = 1'b0;
endcase
casez ({new_n129_, new_n219_})
2'b11 : new_n2651_ = 1'b1;
default : new_n2651_ = 1'b0;
endcase
casez ({v[1], new_n109_})
2'b10 : new_n2652_ = 1'b1;
default : new_n2652_ = 1'b0;
endcase
casez ({new_n162_, new_n220_})
2'b11 : new_n2653_ = 1'b1;
default : new_n2653_ = 1'b0;
endcase
casez ({new_n96_, new_n220_})
2'b11 : new_n2654_ = 1'b1;
default : new_n2654_ = 1'b0;
endcase
casez ({new_n162_, new_n222_})
2'b11 : new_n2655_ = 1'b1;
default : new_n2655_ = 1'b0;
endcase
casez ({new_n221_, new_n223_})
2'b11 : new_n2656_ = 1'b1;
default : new_n2656_ = 1'b0;
endcase
casez ({new_n173_, new_n223_})
2'b11 : new_n2657_ = 1'b1;
default : new_n2657_ = 1'b0;
endcase
casez ({new_n209_, new_n223_})
2'b11 : new_n2658_ = 1'b1;
default : new_n2658_ = 1'b0;
endcase
casez ({new_n144_, new_n223_})
2'b11 : new_n2659_ = 1'b1;
default : new_n2659_ = 1'b0;
endcase
casez ({new_n176_, new_n417_})
2'b11 : new_n2660_ = 1'b1;
default : new_n2660_ = 1'b0;
endcase
casez ({new_n201_, new_n417_})
2'b11 : new_n2661_ = 1'b1;
default : new_n2661_ = 1'b0;
endcase
casez ({new_n196_, new_n417_})
2'b11 : new_n2662_ = 1'b1;
default : new_n2662_ = 1'b0;
endcase
casez ({new_n151_, new_n417_})
2'b11 : new_n2663_ = 1'b1;
default : new_n2663_ = 1'b0;
endcase
casez ({new_n153_, new_n229_})
2'b11 : new_n2664_ = 1'b1;
default : new_n2664_ = 1'b0;
endcase
casez ({new_n151_, new_n432_})
2'b11 : new_n2665_ = 1'b1;
default : new_n2665_ = 1'b0;
endcase
casez ({new_n145_, new_n230_})
2'b11 : new_n2666_ = 1'b1;
default : new_n2666_ = 1'b0;
endcase
casez ({new_n115_, new_n433_})
2'b11 : new_n2667_ = 1'b1;
default : new_n2667_ = 1'b0;
endcase
casez ({new_n82_, new_n237_})
2'b11 : new_n2668_ = 1'b1;
default : new_n2668_ = 1'b0;
endcase
casez ({new_n198_, new_n238_})
2'b11 : new_n2669_ = 1'b1;
default : new_n2669_ = 1'b0;
endcase
casez ({new_n190_, new_n238_})
2'b11 : new_n2670_ = 1'b1;
default : new_n2670_ = 1'b0;
endcase
casez ({new_n170_, new_n241_})
2'b11 : new_n2671_ = 1'b1;
default : new_n2671_ = 1'b0;
endcase
casez ({new_n148_, new_n242_})
2'b11 : new_n2672_ = 1'b1;
default : new_n2672_ = 1'b0;
endcase
casez ({new_n219_, new_n244_})
2'b11 : new_n2673_ = 1'b1;
default : new_n2673_ = 1'b0;
endcase
casez ({new_n137_, new_n469_})
2'b11 : new_n2674_ = 1'b1;
default : new_n2674_ = 1'b0;
endcase
casez ({new_n178_, new_n249_})
2'b11 : new_n2675_ = 1'b1;
default : new_n2675_ = 1'b0;
endcase
casez ({v[1], new_n247_})
2'b01 : new_n2676_ = 1'b1;
default : new_n2676_ = 1'b0;
endcase
casez ({new_n96_, new_n247_})
2'b11 : new_n2677_ = 1'b1;
default : new_n2677_ = 1'b0;
endcase
casez ({y[2], new_n255_})
2'b01 : new_n2678_ = 1'b1;
default : new_n2678_ = 1'b0;
endcase
casez ({new_n123_, new_n142_})
2'b11 : new_n2679_ = 1'b1;
default : new_n2679_ = 1'b0;
endcase
casez ({new_n140_, new_n257_})
2'b11 : new_n2680_ = 1'b1;
default : new_n2680_ = 1'b0;
endcase
casez ({new_n139_, new_n258_})
2'b11 : new_n2681_ = 1'b1;
default : new_n2681_ = 1'b0;
endcase
casez ({new_n118_, new_n258_})
2'b11 : new_n2682_ = 1'b1;
default : new_n2682_ = 1'b0;
endcase
casez ({new_n118_, new_n144_})
2'b11 : new_n2683_ = 1'b1;
default : new_n2683_ = 1'b0;
endcase
casez ({new_n118_, new_n145_})
2'b11 : new_n2684_ = 1'b1;
default : new_n2684_ = 1'b0;
endcase
casez ({y[2], new_n261_})
2'b01 : new_n2685_ = 1'b1;
default : new_n2685_ = 1'b0;
endcase
casez ({new_n133_, new_n146_})
2'b11 : new_n2686_ = 1'b1;
default : new_n2686_ = 1'b0;
endcase
casez ({new_n192_, new_n264_})
2'b11 : new_n2687_ = 1'b1;
default : new_n2687_ = 1'b0;
endcase
casez ({y[2], new_n266_})
2'b01 : new_n2688_ = 1'b1;
default : new_n2688_ = 1'b0;
endcase
casez ({new_n96_, new_n152_})
2'b11 : new_n2689_ = 1'b1;
default : new_n2689_ = 1'b0;
endcase
casez ({new_n144_, new_n153_})
2'b11 : new_n2690_ = 1'b1;
default : new_n2690_ = 1'b0;
endcase
casez ({new_n123_, new_n273_})
2'b11 : new_n2691_ = 1'b1;
default : new_n2691_ = 1'b0;
endcase
casez ({new_n88_, new_n156_})
2'b11 : new_n2692_ = 1'b1;
default : new_n2692_ = 1'b0;
endcase
casez ({new_n159_, new_n274_})
2'b11 : new_n2693_ = 1'b1;
default : new_n2693_ = 1'b0;
endcase
casez ({new_n258_, new_n275_})
2'b11 : new_n2694_ = 1'b1;
default : new_n2694_ = 1'b0;
endcase
casez ({u[2], new_n160_})
2'b01 : new_n2695_ = 1'b1;
default : new_n2695_ = 1'b0;
endcase
casez ({new_n118_, new_n160_})
2'b11 : new_n2696_ = 1'b1;
default : new_n2696_ = 1'b0;
endcase
casez ({y[2], new_n279_})
2'b11 : new_n2697_ = 1'b1;
default : new_n2697_ = 1'b0;
endcase
casez ({new_n150_, new_n161_})
2'b11 : new_n2698_ = 1'b1;
default : new_n2698_ = 1'b0;
endcase
casez ({new_n118_, new_n281_})
2'b11 : new_n2699_ = 1'b1;
default : new_n2699_ = 1'b0;
endcase
casez ({x[2], new_n162_})
2'b01 : new_n2700_ = 1'b1;
default : new_n2700_ = 1'b0;
endcase
casez ({new_n137_, new_n162_})
2'b11 : new_n2701_ = 1'b1;
default : new_n2701_ = 1'b0;
endcase
casez ({new_n139_, new_n161_})
2'b11 : new_n2702_ = 1'b1;
default : new_n2702_ = 1'b0;
endcase
casez ({new_n201_, new_n287_})
2'b11 : new_n2703_ = 1'b1;
default : new_n2703_ = 1'b0;
endcase
casez ({new_n139_, new_n167_})
2'b11 : new_n2704_ = 1'b1;
default : new_n2704_ = 1'b0;
endcase
casez ({new_n123_, new_n167_})
2'b11 : new_n2705_ = 1'b1;
default : new_n2705_ = 1'b0;
endcase
casez ({new_n140_, new_n167_})
2'b11 : new_n2706_ = 1'b1;
default : new_n2706_ = 1'b0;
endcase
casez ({new_n93_, new_n170_})
2'b11 : new_n2707_ = 1'b1;
default : new_n2707_ = 1'b0;
endcase
casez ({new_n159_, new_n299_})
2'b11 : new_n2708_ = 1'b1;
default : new_n2708_ = 1'b0;
endcase
casez ({new_n153_, new_n173_})
2'b11 : new_n2709_ = 1'b1;
default : new_n2709_ = 1'b0;
endcase
casez ({new_n115_, new_n173_})
2'b11 : new_n2710_ = 1'b1;
default : new_n2710_ = 1'b0;
endcase
casez ({new_n118_, new_n176_})
2'b11 : new_n2711_ = 1'b1;
default : new_n2711_ = 1'b0;
endcase
casez ({u[2], new_n177_})
2'b01 : new_n2712_ = 1'b1;
default : new_n2712_ = 1'b0;
endcase
casez ({new_n115_, new_n177_})
2'b11 : new_n2713_ = 1'b1;
default : new_n2713_ = 1'b0;
endcase
casez ({new_n79_, new_n178_})
2'b11 : new_n2714_ = 1'b1;
default : new_n2714_ = 1'b0;
endcase
casez ({new_n118_, new_n178_})
2'b11 : new_n2715_ = 1'b1;
default : new_n2715_ = 1'b0;
endcase
casez ({new_n92_, new_n180_})
2'b11 : new_n2716_ = 1'b1;
default : new_n2716_ = 1'b0;
endcase
casez ({new_n94_, new_n183_})
2'b11 : new_n2717_ = 1'b1;
default : new_n2717_ = 1'b0;
endcase
casez ({new_n229_, new_n328_})
2'b11 : new_n2718_ = 1'b1;
default : new_n2718_ = 1'b0;
endcase
casez ({new_n218_, new_n328_})
2'b11 : new_n2719_ = 1'b1;
default : new_n2719_ = 1'b0;
endcase
casez ({new_n153_, new_n190_})
2'b11 : new_n2720_ = 1'b1;
default : new_n2720_ = 1'b0;
endcase
casez ({new_n142_, new_n189_})
2'b11 : new_n2721_ = 1'b1;
default : new_n2721_ = 1'b0;
endcase
casez ({new_n166_, new_n194_})
2'b11 : new_n2722_ = 1'b1;
default : new_n2722_ = 1'b0;
endcase
casez ({new_n127_, new_n199_})
2'b11 : new_n2723_ = 1'b1;
default : new_n2723_ = 1'b0;
endcase
casez ({new_n94_, new_n343_})
2'b11 : new_n2724_ = 1'b1;
default : new_n2724_ = 1'b0;
endcase
casez ({new_n83_, new_n199_})
2'b11 : new_n2725_ = 1'b1;
default : new_n2725_ = 1'b0;
endcase
casez ({x[1], new_n201_})
2'b11 : new_n2726_ = 1'b1;
default : new_n2726_ = 1'b0;
endcase
casez ({new_n159_, new_n358_})
2'b11 : new_n2727_ = 1'b1;
default : new_n2727_ = 1'b0;
endcase
casez ({new_n144_, new_n363_})
2'b11 : new_n2728_ = 1'b1;
default : new_n2728_ = 1'b0;
endcase
casez ({new_n184_, new_n207_})
2'b11 : new_n2729_ = 1'b1;
default : new_n2729_ = 1'b0;
endcase
casez ({new_n133_, new_n991_})
2'b11 : new_n2730_ = 1'b1;
default : new_n2730_ = 1'b0;
endcase
casez ({new_n103_, new_n209_})
2'b11 : new_n2731_ = 1'b1;
default : new_n2731_ = 1'b0;
endcase
casez ({u[1], new_n211_})
2'b11 : new_n2732_ = 1'b1;
default : new_n2732_ = 1'b0;
endcase
casez ({new_n123_, new_n212_})
2'b11 : new_n2733_ = 1'b1;
default : new_n2733_ = 1'b0;
endcase
casez ({new_n187_, new_n214_})
2'b11 : new_n2734_ = 1'b1;
default : new_n2734_ = 1'b0;
endcase
casez ({new_n209_, new_n215_})
2'b11 : new_n2735_ = 1'b1;
default : new_n2735_ = 1'b0;
endcase
casez ({new_n198_, new_n215_})
2'b11 : new_n2736_ = 1'b1;
default : new_n2736_ = 1'b0;
endcase
casez ({new_n154_, new_n217_})
2'b11 : new_n2737_ = 1'b1;
default : new_n2737_ = 1'b0;
endcase
casez ({new_n85_, new_n219_})
2'b11 : new_n2738_ = 1'b1;
default : new_n2738_ = 1'b0;
endcase
casez ({u[1], new_n219_})
2'b01 : new_n2739_ = 1'b1;
default : new_n2739_ = 1'b0;
endcase
casez ({new_n154_, new_n220_})
2'b11 : new_n2740_ = 1'b1;
default : new_n2740_ = 1'b0;
endcase
casez ({v[1], new_n221_})
2'b01 : new_n2741_ = 1'b1;
default : new_n2741_ = 1'b0;
endcase
casez ({new_n98_, new_n221_})
2'b11 : new_n2742_ = 1'b1;
default : new_n2742_ = 1'b0;
endcase
casez ({u[0], new_n221_})
2'b11 : new_n2743_ = 1'b1;
default : new_n2743_ = 1'b0;
endcase
casez ({new_n198_, new_n229_})
2'b11 : new_n2744_ = 1'b1;
default : new_n2744_ = 1'b0;
endcase
casez ({new_n142_, new_n229_})
2'b11 : new_n2745_ = 1'b1;
default : new_n2745_ = 1'b0;
endcase
casez ({new_n183_, new_n241_})
2'b11 : new_n2746_ = 1'b1;
default : new_n2746_ = 1'b0;
endcase
casez ({u[1], new_n131_})
2'b11 : new_n2747_ = 1'b1;
default : new_n2747_ = 1'b0;
endcase
casez ({new_n89_, new_n243_})
2'b11 : new_n2748_ = 1'b1;
default : new_n2748_ = 1'b0;
endcase
casez ({new_n88_, new_n243_})
2'b11 : new_n2749_ = 1'b1;
default : new_n2749_ = 1'b0;
endcase
casez ({new_n155_, new_n249_})
2'b11 : new_n2750_ = 1'b1;
default : new_n2750_ = 1'b0;
endcase
casez ({new_n187_, new_n249_})
2'b11 : new_n2751_ = 1'b1;
default : new_n2751_ = 1'b0;
endcase
casez ({new_n103_, new_n250_})
2'b11 : new_n2752_ = 1'b1;
default : new_n2752_ = 1'b0;
endcase
casez ({new_n123_, new_n139_})
2'b11 : new_n2753_ = 1'b1;
default : new_n2753_ = 1'b0;
endcase
casez ({new_n97_, new_n144_})
2'b11 : new_n2754_ = 1'b1;
default : new_n2754_ = 1'b0;
endcase
casez ({x[2], new_n150_})
2'b11 : new_n2755_ = 1'b1;
default : new_n2755_ = 1'b0;
endcase
casez ({new_n104_, new_n150_})
2'b11 : new_n2756_ = 1'b1;
default : new_n2756_ = 1'b0;
endcase
casez ({y[2], new_n155_})
2'b01 : new_n2757_ = 1'b1;
default : new_n2757_ = 1'b0;
endcase
casez ({new_n95_, new_n160_})
2'b11 : new_n2758_ = 1'b1;
default : new_n2758_ = 1'b0;
endcase
casez ({new_n80_, new_n166_})
2'b11 : new_n2759_ = 1'b1;
default : new_n2759_ = 1'b0;
endcase
casez ({u[2], new_n176_})
2'b01 : new_n2760_ = 1'b1;
default : new_n2760_ = 1'b0;
endcase
casez ({new_n83_, new_n182_})
2'b11 : new_n2761_ = 1'b1;
default : new_n2761_ = 1'b0;
endcase
casez ({u[2], new_n183_})
2'b11 : new_n2762_ = 1'b1;
default : new_n2762_ = 1'b0;
endcase
casez ({new_n80_, new_n184_})
2'b11 : new_n2763_ = 1'b1;
default : new_n2763_ = 1'b0;
endcase
casez ({u[2], new_n200_})
2'b11 : new_n2764_ = 1'b1;
default : new_n2764_ = 1'b0;
endcase
casez ({new_n92_, new_n204_})
2'b11 : new_n2765_ = 1'b1;
default : new_n2765_ = 1'b0;
endcase
casez ({new_n88_, new_n115_})
2'b11 : new_n2766_ = 1'b1;
default : new_n2766_ = 1'b0;
endcase
casez ({u[1], new_n118_})
2'b11 : new_n2767_ = 1'b1;
default : new_n2767_ = 1'b0;
endcase
casez ({new_n103_, new_n118_})
2'b11 : new_n2768_ = 1'b1;
default : new_n2768_ = 1'b0;
endcase
casez ({new_n104_, new_n118_})
2'b11 : new_n2769_ = 1'b1;
default : new_n2769_ = 1'b0;
endcase
casez ({new_n80_, new_n120_})
2'b11 : new_n2770_ = 1'b1;
default : new_n2770_ = 1'b0;
endcase
casez ({y[2], new_n123_})
2'b01 : new_n2771_ = 1'b1;
default : new_n2771_ = 1'b0;
endcase
casez ({new_n79_, new_n123_})
2'b11 : new_n2772_ = 1'b1;
default : new_n2772_ = 1'b0;
endcase
casez ({new_n89_, new_n126_})
2'b11 : new_n2773_ = 1'b1;
default : new_n2773_ = 1'b0;
endcase
casez ({new_n96_, new_n126_})
2'b11 : new_n2774_ = 1'b1;
default : new_n2774_ = 1'b0;
endcase
casez ({new_n92_, new_n128_})
2'b11 : new_n2775_ = 1'b1;
default : new_n2775_ = 1'b0;
endcase
casez ({new_n89_, new_n131_})
2'b11 : new_n2776_ = 1'b1;
default : new_n2776_ = 1'b0;
endcase
casez ({new_n84_, new_n137_})
2'b11 : new_n2777_ = 1'b1;
default : new_n2777_ = 1'b0;
endcase
casez ({new_n81_, new_n115_})
2'b11 : new_n2778_ = 1'b1;
default : new_n2778_ = 1'b0;
endcase
casez ({new_n85_, new_n115_})
2'b11 : new_n2779_ = 1'b1;
default : new_n2779_ = 1'b0;
endcase
casez ({v[1], new_n127_})
2'b01 : new_n2780_ = 1'b1;
default : new_n2780_ = 1'b0;
endcase
casez ({new_n96_, new_n430_, new_n101_, new_n604_})
4'b11?? : new_n2781_ = 1'b1;
4'b??11 : new_n2781_ = 1'b1;
default : new_n2781_ = 1'b0;
endcase
casez ({new_n228_, new_n360_})
2'b00 : new_n2782_ = 1'b1;
default : new_n2782_ = 1'b0;
endcase
casez ({new_n311_, new_n361_})
2'b00 : new_n2783_ = 1'b1;
default : new_n2783_ = 1'b0;
endcase
casez ({new_n173_, new_n672_})
2'b00 : new_n2784_ = 1'b1;
default : new_n2784_ = 1'b0;
endcase
casez ({new_n274_, new_n388_})
2'b00 : new_n2785_ = 1'b1;
default : new_n2785_ = 1'b0;
endcase
casez ({new_n273_, new_n430_})
2'b00 : new_n2786_ = 1'b1;
default : new_n2786_ = 1'b0;
endcase
casez ({new_n103_, new_n505_})
2'b11 : new_n2787_ = 1'b1;
default : new_n2787_ = 1'b0;
endcase
casez ({new_n91_, new_n526_})
2'b11 : new_n2788_ = 1'b1;
default : new_n2788_ = 1'b0;
endcase
casez ({new_n85_, new_n541_})
2'b11 : new_n2789_ = 1'b1;
default : new_n2789_ = 1'b0;
endcase
casez ({v[0], new_n542_})
2'b11 : new_n2790_ = 1'b1;
default : new_n2790_ = 1'b0;
endcase
casez ({new_n81_, new_n555_})
2'b01 : new_n2791_ = 1'b1;
default : new_n2791_ = 1'b0;
endcase
casez ({x[2], new_n290_})
2'b11 : new_n2792_ = 1'b1;
default : new_n2792_ = 1'b0;
endcase
casez ({y[1], new_n308_})
2'b11 : new_n2793_ = 1'b1;
default : new_n2793_ = 1'b0;
endcase
casez ({new_n86_, new_n605_})
2'b11 : new_n2794_ = 1'b1;
default : new_n2794_ = 1'b0;
endcase
casez ({x[0], new_n181_})
2'b10 : new_n2795_ = 1'b1;
default : new_n2795_ = 1'b0;
endcase
casez ({y[1], new_n329_})
2'b11 : new_n2796_ = 1'b1;
default : new_n2796_ = 1'b0;
endcase
casez ({x[0], new_n671_})
2'b11 : new_n2797_ = 1'b1;
default : new_n2797_ = 1'b0;
endcase
casez ({new_n84_, new_n678_})
2'b01 : new_n2798_ = 1'b1;
default : new_n2798_ = 1'b0;
endcase
casez ({y[1], new_n395_})
2'b11 : new_n2799_ = 1'b1;
default : new_n2799_ = 1'b0;
endcase
casez ({new_n105_, new_n395_})
2'b11 : new_n2800_ = 1'b1;
default : new_n2800_ = 1'b0;
endcase
casez ({new_n120_, new_n397_})
2'b11 : new_n2801_ = 1'b1;
default : new_n2801_ = 1'b0;
endcase
casez ({y[0], new_n397_})
2'b11 : new_n2802_ = 1'b1;
default : new_n2802_ = 1'b0;
endcase
casez ({v[0], new_n1045_})
2'b11 : new_n2803_ = 1'b1;
default : new_n2803_ = 1'b0;
endcase
casez ({new_n91_, new_n421_})
2'b11 : new_n2804_ = 1'b1;
default : new_n2804_ = 1'b0;
endcase
casez ({u[2], new_n421_})
2'b11 : new_n2805_ = 1'b1;
default : new_n2805_ = 1'b0;
endcase
casez ({new_n169_, new_n422_})
2'b11 : new_n2806_ = 1'b1;
default : new_n2806_ = 1'b0;
endcase
casez ({v[2], new_n741_})
2'b01 : new_n2807_ = 1'b1;
default : new_n2807_ = 1'b0;
endcase
casez ({y[1], new_n741_})
2'b11 : new_n2808_ = 1'b1;
default : new_n2808_ = 1'b0;
endcase
casez ({new_n80_, new_n745_})
2'b01 : new_n2809_ = 1'b1;
default : new_n2809_ = 1'b0;
endcase
casez ({new_n86_, new_n481_})
2'b11 : new_n2810_ = 1'b1;
default : new_n2810_ = 1'b0;
endcase
casez ({new_n89_, new_n781_})
2'b11 : new_n2811_ = 1'b1;
default : new_n2811_ = 1'b0;
endcase
casez ({new_n107_, new_n259_})
2'b01 : new_n2812_ = 1'b1;
default : new_n2812_ = 1'b0;
endcase
casez ({new_n92_, new_n259_})
2'b11 : new_n2813_ = 1'b1;
default : new_n2813_ = 1'b0;
endcase
casez ({new_n98_, new_n265_})
2'b11 : new_n2814_ = 1'b1;
default : new_n2814_ = 1'b0;
endcase
casez ({y[0], new_n526_})
2'b01 : new_n2815_ = 1'b1;
default : new_n2815_ = 1'b0;
endcase
casez ({u[0], new_n527_})
2'b11 : new_n2816_ = 1'b1;
default : new_n2816_ = 1'b0;
endcase
casez ({new_n114_, new_n156_})
2'b11 : new_n2817_ = 1'b1;
default : new_n2817_ = 1'b0;
endcase
casez ({new_n84_, new_n551_})
2'b11 : new_n2818_ = 1'b1;
default : new_n2818_ = 1'b0;
endcase
casez ({new_n186_, new_n287_})
2'b11 : new_n2819_ = 1'b1;
default : new_n2819_ = 1'b0;
endcase
casez ({v[1], new_n294_})
2'b01 : new_n2820_ = 1'b1;
default : new_n2820_ = 1'b0;
endcase
casez ({new_n77_, new_n308_})
2'b11 : new_n2821_ = 1'b1;
default : new_n2821_ = 1'b0;
endcase
casez ({y[2], new_n603_})
2'b11 : new_n2822_ = 1'b1;
default : new_n2822_ = 1'b0;
endcase
casez ({new_n186_, new_n317_})
2'b11 : new_n2823_ = 1'b1;
default : new_n2823_ = 1'b0;
endcase
casez ({new_n101_, new_n335_})
2'b11 : new_n2824_ = 1'b1;
default : new_n2824_ = 1'b0;
endcase
casez ({new_n88_, new_n340_})
2'b11 : new_n2825_ = 1'b1;
default : new_n2825_ = 1'b0;
endcase
casez ({new_n187_, new_n360_})
2'b11 : new_n2826_ = 1'b1;
default : new_n2826_ = 1'b0;
endcase
casez ({new_n86_, new_n378_})
2'b11 : new_n2827_ = 1'b1;
default : new_n2827_ = 1'b0;
endcase
casez ({new_n171_, new_n211_})
2'b11 : new_n2828_ = 1'b1;
default : new_n2828_ = 1'b0;
endcase
casez ({new_n85_, new_n381_})
2'b11 : new_n2829_ = 1'b1;
default : new_n2829_ = 1'b0;
endcase
casez ({new_n186_, new_n212_})
2'b11 : new_n2830_ = 1'b1;
default : new_n2830_ = 1'b0;
endcase
casez ({u[0], new_n383_})
2'b11 : new_n2831_ = 1'b1;
default : new_n2831_ = 1'b0;
endcase
casez ({x[0], new_n390_})
2'b01 : new_n2832_ = 1'b1;
default : new_n2832_ = 1'b0;
endcase
casez ({new_n100_, new_n397_})
2'b11 : new_n2833_ = 1'b1;
default : new_n2833_ = 1'b0;
endcase
casez ({v[0], new_n408_})
2'b01 : new_n2834_ = 1'b1;
default : new_n2834_ = 1'b0;
endcase
casez ({new_n97_, new_n420_})
2'b11 : new_n2835_ = 1'b1;
default : new_n2835_ = 1'b0;
endcase
casez ({new_n97_, new_n428_})
2'b10 : new_n2836_ = 1'b1;
default : new_n2836_ = 1'b0;
endcase
casez ({new_n96_, new_n435_})
2'b11 : new_n2837_ = 1'b1;
default : new_n2837_ = 1'b0;
endcase
casez ({y[2], new_n439_})
2'b00 : new_n2838_ = 1'b1;
default : new_n2838_ = 1'b0;
endcase
casez ({u[1], new_n719_})
2'b11 : new_n2839_ = 1'b1;
default : new_n2839_ = 1'b0;
endcase
casez ({v[2], new_n449_})
2'b01 : new_n2840_ = 1'b1;
default : new_n2840_ = 1'b0;
endcase
casez ({new_n82_, new_n449_})
2'b01 : new_n2841_ = 1'b1;
default : new_n2841_ = 1'b0;
endcase
casez ({x[1], new_n456_})
2'b11 : new_n2842_ = 1'b1;
default : new_n2842_ = 1'b0;
endcase
casez ({new_n103_, new_n460_})
2'b11 : new_n2843_ = 1'b1;
default : new_n2843_ = 1'b0;
endcase
casez ({new_n137_, new_n1119_})
2'b11 : new_n2844_ = 1'b1;
default : new_n2844_ = 1'b0;
endcase
casez ({new_n112_, new_n250_})
2'b11 : new_n2845_ = 1'b1;
default : new_n2845_ = 1'b0;
endcase
casez ({u[2], new_n259_})
2'b01 : new_n2846_ = 1'b1;
default : new_n2846_ = 1'b0;
endcase
casez ({new_n83_, new_n268_})
2'b11 : new_n2847_ = 1'b1;
default : new_n2847_ = 1'b0;
endcase
casez ({new_n83_, new_n323_})
2'b11 : new_n2848_ = 1'b1;
default : new_n2848_ = 1'b0;
endcase
casez ({new_n79_, new_n545_})
2'b11 : new_n2849_ = 1'b1;
default : new_n2849_ = 1'b0;
endcase
casez ({new_n384_, new_n546_})
2'b00 : new_n2850_ = 1'b1;
default : new_n2850_ = 1'b0;
endcase
casez ({new_n355_, new_n425_})
2'b00 : new_n2851_ = 1'b1;
default : new_n2851_ = 1'b0;
endcase
casez ({new_n144_, new_n1687_, new_n1968_})
3'b11? : new_n2852_ = 1'b1;
3'b??1 : new_n2852_ = 1'b1;
default : new_n2852_ = 1'b0;
endcase
casez ({new_n312_, new_n795_, new_n1977_})
3'b11? : new_n2853_ = 1'b1;
3'b??1 : new_n2853_ = 1'b1;
default : new_n2853_ = 1'b0;
endcase
casez ({new_n322_, new_n703_, new_n1985_})
3'b11? : new_n2854_ = 1'b1;
3'b??1 : new_n2854_ = 1'b1;
default : new_n2854_ = 1'b0;
endcase
casez ({new_n211_, new_n1063_, new_n1989_})
3'b11? : new_n2855_ = 1'b1;
3'b??1 : new_n2855_ = 1'b1;
default : new_n2855_ = 1'b0;
endcase
casez ({new_n335_, new_n990_, new_n2002_})
3'b11? : new_n2856_ = 1'b1;
3'b??1 : new_n2856_ = 1'b1;
default : new_n2856_ = 1'b0;
endcase
casez ({new_n480_, new_n1108_, new_n2007_})
3'b11? : new_n2857_ = 1'b1;
3'b??1 : new_n2857_ = 1'b1;
default : new_n2857_ = 1'b0;
endcase
casez ({v[2], new_n1442_, new_n2016_})
3'b11? : new_n2858_ = 1'b1;
3'b??1 : new_n2858_ = 1'b1;
default : new_n2858_ = 1'b0;
endcase
casez ({new_n342_, new_n463_, new_n2020_})
3'b11? : new_n2859_ = 1'b1;
3'b??1 : new_n2859_ = 1'b1;
default : new_n2859_ = 1'b0;
endcase
casez ({new_n171_, new_n1632_, new_n2021_})
3'b11? : new_n2860_ = 1'b1;
3'b??1 : new_n2860_ = 1'b1;
default : new_n2860_ = 1'b0;
endcase
casez ({new_n239_, new_n1524_, new_n2023_})
3'b11? : new_n2861_ = 1'b1;
3'b??1 : new_n2861_ = 1'b1;
default : new_n2861_ = 1'b0;
endcase
casez ({new_n187_, new_n518_, new_n2030_})
3'b11? : new_n2862_ = 1'b1;
3'b??1 : new_n2862_ = 1'b1;
default : new_n2862_ = 1'b0;
endcase
casez ({new_n390_, new_n982_, new_n2034_})
3'b11? : new_n2863_ = 1'b1;
3'b??1 : new_n2863_ = 1'b1;
default : new_n2863_ = 1'b0;
endcase
casez ({new_n183_, new_n1269_, new_n2042_})
3'b11? : new_n2864_ = 1'b1;
3'b??1 : new_n2864_ = 1'b1;
default : new_n2864_ = 1'b0;
endcase
casez ({new_n194_, new_n1068_, new_n2088_})
3'b11? : new_n2865_ = 1'b1;
3'b??1 : new_n2865_ = 1'b1;
default : new_n2865_ = 1'b0;
endcase
casez ({new_n459_, new_n653_, new_n2100_})
3'b11? : new_n2866_ = 1'b1;
3'b??1 : new_n2866_ = 1'b1;
default : new_n2866_ = 1'b0;
endcase
casez ({new_n249_, new_n2139_, new_n2018_})
3'b11? : new_n2867_ = 1'b1;
3'b??1 : new_n2867_ = 1'b1;
default : new_n2867_ = 1'b0;
endcase
casez ({new_n179_, new_n474_, new_n1128_})
3'b11? : new_n2868_ = 1'b1;
3'b??1 : new_n2868_ = 1'b1;
default : new_n2868_ = 1'b0;
endcase
casez ({new_n79_, new_n485_})
2'b10 : new_n2869_ = 1'b1;
default : new_n2869_ = 1'b0;
endcase
casez ({new_n234_, new_n443_})
2'b11 : new_n2870_ = 1'b1;
default : new_n2870_ = 1'b0;
endcase
casez ({new_n1232_, new_n1233_})
2'b00 : new_n2871_ = 1'b1;
default : new_n2871_ = 1'b0;
endcase
casez ({new_n189_, new_n917_, new_n2173_})
3'b11? : new_n2872_ = 1'b1;
3'b??1 : new_n2872_ = 1'b1;
default : new_n2872_ = 1'b0;
endcase
casez ({new_n157_, new_n587_, new_n2177_})
3'b11? : new_n2873_ = 1'b1;
3'b??1 : new_n2873_ = 1'b1;
default : new_n2873_ = 1'b0;
endcase
casez ({new_n6129_, new_n2192_})
2'b1? : new_n2874_ = 1'b1;
2'b?1 : new_n2874_ = 1'b1;
default : new_n2874_ = 1'b0;
endcase
casez ({new_n299_, new_n2145_, new_n2196_})
3'b11? : new_n2875_ = 1'b1;
3'b??1 : new_n2875_ = 1'b1;
default : new_n2875_ = 1'b0;
endcase
casez ({new_n371_, new_n1688_, new_n2197_})
3'b11? : new_n2876_ = 1'b1;
3'b??1 : new_n2876_ = 1'b1;
default : new_n2876_ = 1'b0;
endcase
casez ({new_n223_, new_n1786_, new_n2204_})
3'b11? : new_n2877_ = 1'b1;
3'b??1 : new_n2877_ = 1'b1;
default : new_n2877_ = 1'b0;
endcase
casez ({new_n238_, new_n1082_, new_n2215_})
3'b10? : new_n2878_ = 1'b1;
3'b??1 : new_n2878_ = 1'b1;
default : new_n2878_ = 1'b0;
endcase
casez ({new_n350_, new_n912_, new_n2218_})
3'b11? : new_n2879_ = 1'b1;
3'b??1 : new_n2879_ = 1'b1;
default : new_n2879_ = 1'b0;
endcase
casez ({new_n236_, new_n1053_, new_n2239_})
3'b10? : new_n2880_ = 1'b1;
3'b??1 : new_n2880_ = 1'b1;
default : new_n2880_ = 1'b0;
endcase
casez ({new_n122_, new_n1450_, new_n2242_})
3'b11? : new_n2881_ = 1'b1;
3'b??1 : new_n2881_ = 1'b1;
default : new_n2881_ = 1'b0;
endcase
casez ({new_n385_, new_n1140_, new_n2268_})
3'b11? : new_n2882_ = 1'b1;
3'b??1 : new_n2882_ = 1'b1;
default : new_n2882_ = 1'b0;
endcase
casez ({new_n228_, new_n645_, new_n2270_})
3'b11? : new_n2883_ = 1'b1;
3'b??1 : new_n2883_ = 1'b1;
default : new_n2883_ = 1'b0;
endcase
casez ({new_n132_, new_n1123_, new_n2289_})
3'b11? : new_n2884_ = 1'b1;
3'b??1 : new_n2884_ = 1'b1;
default : new_n2884_ = 1'b0;
endcase
casez ({new_n208_, new_n1072_, new_n2296_})
3'b11? : new_n2885_ = 1'b1;
3'b??1 : new_n2885_ = 1'b1;
default : new_n2885_ = 1'b0;
endcase
casez ({new_n307_, new_n546_, new_n2310_})
3'b11? : new_n2886_ = 1'b1;
3'b??1 : new_n2886_ = 1'b1;
default : new_n2886_ = 1'b0;
endcase
casez ({new_n334_, new_n1087_, new_n2329_})
3'b11? : new_n2887_ = 1'b1;
3'b??1 : new_n2887_ = 1'b1;
default : new_n2887_ = 1'b0;
endcase
casez ({new_n550_, new_n1762_, new_n2332_})
3'b00? : new_n2888_ = 1'b1;
3'b??1 : new_n2888_ = 1'b1;
default : new_n2888_ = 1'b0;
endcase
casez ({new_n731_, new_n1234_})
2'b00 : new_n2889_ = 1'b1;
default : new_n2889_ = 1'b0;
endcase
casez ({new_n1240_, new_n1779_})
2'b00 : new_n2890_ = 1'b1;
default : new_n2890_ = 1'b0;
endcase
casez ({new_n169_, new_n1537_, new_n1995_})
3'b11? : new_n2891_ = 1'b1;
3'b??1 : new_n2891_ = 1'b1;
default : new_n2891_ = 1'b0;
endcase
casez ({new_n263_, new_n646_, new_n1246_})
3'b11? : new_n2892_ = 1'b1;
3'b??1 : new_n2892_ = 1'b1;
default : new_n2892_ = 1'b0;
endcase
casez ({new_n100_, new_n1006_, new_n1251_})
3'b11? : new_n2893_ = 1'b1;
3'b??1 : new_n2893_ = 1'b1;
default : new_n2893_ = 1'b0;
endcase
casez ({new_n224_, new_n849_, new_n2341_})
3'b11? : new_n2894_ = 1'b1;
3'b??1 : new_n2894_ = 1'b1;
default : new_n2894_ = 1'b0;
endcase
casez ({new_n90_, new_n466_, new_n2350_})
3'b11? : new_n2895_ = 1'b1;
3'b??1 : new_n2895_ = 1'b1;
default : new_n2895_ = 1'b0;
endcase
casez ({new_n401_, new_n642_, new_n2353_})
3'b11? : new_n2896_ = 1'b1;
3'b??1 : new_n2896_ = 1'b1;
default : new_n2896_ = 1'b0;
endcase
casez ({new_n241_, new_n951_, new_n2359_})
3'b11? : new_n2897_ = 1'b1;
3'b??1 : new_n2897_ = 1'b1;
default : new_n2897_ = 1'b0;
endcase
casez ({new_n118_, new_n1068_, new_n2362_})
3'b11? : new_n2898_ = 1'b1;
3'b??1 : new_n2898_ = 1'b1;
default : new_n2898_ = 1'b0;
endcase
casez ({new_n268_, new_n446_, new_n2398_})
3'b11? : new_n2899_ = 1'b1;
3'b??1 : new_n2899_ = 1'b1;
default : new_n2899_ = 1'b0;
endcase
casez ({new_n386_, new_n1887_, new_n2407_})
3'b11? : new_n2900_ = 1'b1;
3'b??1 : new_n2900_ = 1'b1;
default : new_n2900_ = 1'b0;
endcase
casez ({new_n85_, new_n1509_, new_n2424_})
3'b11? : new_n2901_ = 1'b1;
3'b??1 : new_n2901_ = 1'b1;
default : new_n2901_ = 1'b0;
endcase
casez ({new_n104_, new_n1789_, new_n2391_})
3'b11? : new_n2902_ = 1'b1;
3'b??1 : new_n2902_ = 1'b1;
default : new_n2902_ = 1'b0;
endcase
casez ({new_n137_, new_n466_, new_n2439_})
3'b11? : new_n2903_ = 1'b1;
3'b??1 : new_n2903_ = 1'b1;
default : new_n2903_ = 1'b0;
endcase
casez ({new_n179_, new_n1563_, new_n2444_})
3'b11? : new_n2904_ = 1'b1;
3'b??1 : new_n2904_ = 1'b1;
default : new_n2904_ = 1'b0;
endcase
casez ({new_n427_, new_n614_, new_n2452_})
3'b11? : new_n2905_ = 1'b1;
3'b??1 : new_n2905_ = 1'b1;
default : new_n2905_ = 1'b0;
endcase
casez ({new_n192_, new_n514_, new_n2472_})
3'b11? : new_n2906_ = 1'b1;
3'b??1 : new_n2906_ = 1'b1;
default : new_n2906_ = 1'b0;
endcase
casez ({new_n398_, new_n1740_, new_n2476_})
3'b11? : new_n2907_ = 1'b1;
3'b??1 : new_n2907_ = 1'b1;
default : new_n2907_ = 1'b0;
endcase
casez ({new_n448_, new_n810_, new_n1493_})
3'b11? : new_n2908_ = 1'b1;
3'b??1 : new_n2908_ = 1'b1;
default : new_n2908_ = 1'b0;
endcase
casez ({new_n217_, new_n546_, new_n1791_})
3'b11? : new_n2909_ = 1'b1;
3'b??1 : new_n2909_ = 1'b1;
default : new_n2909_ = 1'b0;
endcase
casez ({new_n183_, new_n697_, new_n1792_})
3'b11? : new_n2910_ = 1'b1;
3'b??1 : new_n2910_ = 1'b1;
default : new_n2910_ = 1'b0;
endcase
casez ({new_n97_, new_n1795_, new_n2174_})
3'b11? : new_n2911_ = 1'b1;
3'b??1 : new_n2911_ = 1'b1;
default : new_n2911_ = 1'b0;
endcase
casez ({x[1], y[2]})
2'b01 : new_n2912_ = 1'b1;
default : new_n2912_ = 1'b0;
endcase
casez ({y[0], y[1]})
2'b10 : new_n2913_ = 1'b1;
default : new_n2913_ = 1'b0;
endcase
casez ({x[1], u[0]})
2'b01 : new_n2914_ = 1'b1;
default : new_n2914_ = 1'b0;
endcase
casez ({x[1], x[2]})
2'b00 : new_n2915_ = 1'b1;
default : new_n2915_ = 1'b0;
endcase
casez ({y[0], y[1]})
2'b01 : new_n2916_ = 1'b1;
default : new_n2916_ = 1'b0;
endcase
casez ({u[0], u[2]})
2'b00 : new_n2917_ = 1'b1;
default : new_n2917_ = 1'b0;
endcase
casez ({new_n79_, new_n85_})
2'b00 : new_n2918_ = 1'b1;
default : new_n2918_ = 1'b0;
endcase
casez ({x[1], new_n86_, x[2], u[2]})
4'b01?? : new_n2919_ = 1'b1;
4'b??01 : new_n2919_ = 1'b1;
default : new_n2919_ = 1'b0;
endcase
casez ({new_n2961_, new_n234_})
2'b1? : new_n2920_ = 1'b1;
2'b?1 : new_n2920_ = 1'b1;
default : new_n2920_ = 1'b0;
endcase
casez ({new_n2974_, new_n2959_})
2'b1? : new_n2921_ = 1'b1;
2'b?1 : new_n2921_ = 1'b1;
default : new_n2921_ = 1'b0;
endcase
casez ({new_n79_, new_n104_, new_n92_, new_n278_})
4'b01?? : new_n2922_ = 1'b1;
4'b??01 : new_n2922_ = 1'b1;
default : new_n2922_ = 1'b0;
endcase
casez ({new_n2978_, new_n2496_})
2'b1? : new_n2923_ = 1'b1;
2'b?1 : new_n2923_ = 1'b1;
default : new_n2923_ = 1'b0;
endcase
casez ({new_n2967_, new_n437_})
2'b1? : new_n2924_ = 1'b1;
2'b?1 : new_n2924_ = 1'b1;
default : new_n2924_ = 1'b0;
endcase
casez ({new_n86_, new_n1796_, new_n104_, new_n1257_})
4'b11?? : new_n2925_ = 1'b1;
4'b??11 : new_n2925_ = 1'b1;
default : new_n2925_ = 1'b0;
endcase
casez ({new_n97_, new_n257_})
2'b00 : new_n2926_ = 1'b1;
default : new_n2926_ = 1'b0;
endcase
casez ({new_n487_, new_n1539_})
2'b00 : new_n2927_ = 1'b1;
default : new_n2927_ = 1'b0;
endcase
casez ({new_n98_, new_n444_})
2'b00 : new_n2928_ = 1'b1;
default : new_n2928_ = 1'b0;
endcase
casez ({new_n89_, new_n346_})
2'b00 : new_n2929_ = 1'b1;
default : new_n2929_ = 1'b0;
endcase
casez ({new_n88_, new_n224_})
2'b00 : new_n2930_ = 1'b1;
default : new_n2930_ = 1'b0;
endcase
casez ({new_n224_, new_n242_})
2'b00 : new_n2931_ = 1'b1;
default : new_n2931_ = 1'b0;
endcase
casez ({v[1], new_n93_})
2'b11 : new_n2932_ = 1'b1;
default : new_n2932_ = 1'b0;
endcase
casez ({new_n81_, new_n91_})
2'b01 : new_n2933_ = 1'b1;
default : new_n2933_ = 1'b0;
endcase
casez ({x[2], new_n92_})
2'b10 : new_n2934_ = 1'b1;
default : new_n2934_ = 1'b0;
endcase
casez ({v[2], new_n97_})
2'b01 : new_n2935_ = 1'b1;
default : new_n2935_ = 1'b0;
endcase
casez ({v[1], new_n79_})
2'b00 : new_n2936_ = 1'b1;
default : new_n2936_ = 1'b0;
endcase
casez ({y[2], new_n79_})
2'b10 : new_n2937_ = 1'b1;
default : new_n2937_ = 1'b0;
endcase
casez ({new_n81_, new_n98_})
2'b01 : new_n2938_ = 1'b1;
default : new_n2938_ = 1'b0;
endcase
casez ({v[1], new_n80_})
2'b00 : new_n2939_ = 1'b1;
default : new_n2939_ = 1'b0;
endcase
casez ({v[2], new_n101_})
2'b01 : new_n2940_ = 1'b1;
default : new_n2940_ = 1'b0;
endcase
casez ({x[1], new_n104_})
2'b01 : new_n2941_ = 1'b1;
default : new_n2941_ = 1'b0;
endcase
casez ({new_n84_, new_n104_})
2'b11 : new_n2942_ = 1'b1;
default : new_n2942_ = 1'b0;
endcase
casez ({new_n92_, new_n104_})
2'b11 : new_n2943_ = 1'b1;
default : new_n2943_ = 1'b0;
endcase
casez ({v[0], new_n82_})
2'b10 : new_n2944_ = 1'b1;
default : new_n2944_ = 1'b0;
endcase
casez ({v[0], new_n257_})
2'b01 : new_n2945_ = 1'b1;
default : new_n2945_ = 1'b0;
endcase
casez ({u[1], new_n96_})
2'b00 : new_n2946_ = 1'b1;
default : new_n2946_ = 1'b0;
endcase
casez ({new_n93_, new_n346_})
2'b11 : new_n2947_ = 1'b1;
default : new_n2947_ = 1'b0;
endcase
casez ({new_n85_, new_n101_})
2'b01 : new_n2948_ = 1'b1;
default : new_n2948_ = 1'b0;
endcase
casez ({new_n80_, new_n103_})
2'b01 : new_n2949_ = 1'b1;
default : new_n2949_ = 1'b0;
endcase
casez ({u[0], new_n104_})
2'b10 : new_n2950_ = 1'b1;
default : new_n2950_ = 1'b0;
endcase
casez ({u[0], new_n104_})
2'b01 : new_n2951_ = 1'b1;
default : new_n2951_ = 1'b0;
endcase
casez ({u[2], new_n230_})
2'b01 : new_n2952_ = 1'b1;
default : new_n2952_ = 1'b0;
endcase
casez ({new_n83_, new_n234_})
2'b11 : new_n2953_ = 1'b1;
default : new_n2953_ = 1'b0;
endcase
casez ({new_n97_, new_n234_})
2'b11 : new_n2954_ = 1'b1;
default : new_n2954_ = 1'b0;
endcase
casez ({u[0], new_n85_})
2'b10 : new_n2955_ = 1'b1;
default : new_n2955_ = 1'b0;
endcase
casez ({x[1], new_n242_})
2'b11 : new_n2956_ = 1'b1;
default : new_n2956_ = 1'b0;
endcase
casez ({new_n93_, new_n242_})
2'b11 : new_n2957_ = 1'b1;
default : new_n2957_ = 1'b0;
endcase
casez ({new_n98_, new_n487_})
2'b11 : new_n2958_ = 1'b1;
default : new_n2958_ = 1'b0;
endcase
casez ({new_n98_, new_n486_})
2'b11 : new_n2959_ = 1'b1;
default : new_n2959_ = 1'b0;
endcase
casez ({new_n81_, new_n91_})
2'b10 : new_n2960_ = 1'b1;
default : new_n2960_ = 1'b0;
endcase
casez ({x[1], new_n284_})
2'b01 : new_n2961_ = 1'b1;
default : new_n2961_ = 1'b0;
endcase
casez ({new_n91_, new_n94_})
2'b10 : new_n2962_ = 1'b1;
default : new_n2962_ = 1'b0;
endcase
casez ({new_n90_, new_n94_})
2'b10 : new_n2963_ = 1'b1;
default : new_n2963_ = 1'b0;
endcase
casez ({new_n90_, new_n95_})
2'b01 : new_n2964_ = 1'b1;
default : new_n2964_ = 1'b0;
endcase
casez ({u[1], new_n923_})
2'b01 : new_n2965_ = 1'b1;
default : new_n2965_ = 1'b0;
endcase
casez ({new_n85_, new_n923_})
2'b11 : new_n2966_ = 1'b1;
default : new_n2966_ = 1'b0;
endcase
casez ({y[1], new_n99_})
2'b11 : new_n2967_ = 1'b1;
default : new_n2967_ = 1'b0;
endcase
casez ({new_n86_, new_n101_})
2'b10 : new_n2968_ = 1'b1;
default : new_n2968_ = 1'b0;
endcase
casez ({new_n79_, new_n230_})
2'b01 : new_n2969_ = 1'b1;
default : new_n2969_ = 1'b0;
endcase
casez ({u[1], new_n728_})
2'b01 : new_n2970_ = 1'b1;
default : new_n2970_ = 1'b0;
endcase
casez ({y[1], new_n1090_})
2'b11 : new_n2971_ = 1'b1;
default : new_n2971_ = 1'b0;
endcase
casez ({new_n89_, new_n92_})
2'b11 : new_n2972_ = 1'b1;
default : new_n2972_ = 1'b0;
endcase
casez ({u[1], new_n93_})
2'b01 : new_n2973_ = 1'b1;
default : new_n2973_ = 1'b0;
endcase
casez ({v[1], new_n95_})
2'b01 : new_n2974_ = 1'b1;
default : new_n2974_ = 1'b0;
endcase
casez ({y[0], new_n97_})
2'b01 : new_n2975_ = 1'b1;
default : new_n2975_ = 1'b0;
endcase
casez ({v[1], new_n100_})
2'b01 : new_n2976_ = 1'b1;
default : new_n2976_ = 1'b0;
endcase
casez ({x[1], new_n101_})
2'b11 : new_n2977_ = 1'b1;
default : new_n2977_ = 1'b0;
endcase
casez ({x[1], new_n85_})
2'b11 : new_n2978_ = 1'b1;
default : new_n2978_ = 1'b0;
endcase
casez ({new_n79_, new_n86_})
2'b11 : new_n2979_ = 1'b1;
default : new_n2979_ = 1'b0;
endcase
casez ({x[2], new_n79_})
2'b11 : new_n2980_ = 1'b1;
default : new_n2980_ = 1'b0;
endcase
casez ({u[1], new_n80_, new_n135_})
3'b11? : new_n2981_ = 1'b1;
3'b??1 : new_n2981_ = 1'b1;
default : new_n2981_ = 1'b0;
endcase
casez ({new_n204_, new_n764_, new_n3393_})
3'b11? : new_n2982_ = 1'b1;
3'b??1 : new_n2982_ = 1'b1;
default : new_n2982_ = 1'b0;
endcase
casez ({new_n187_, new_n251_})
2'b00 : new_n2983_ = 1'b1;
default : new_n2983_ = 1'b0;
endcase
casez ({new_n198_, new_n237_, new_n767_})
3'b11? : new_n2984_ = 1'b1;
3'b??1 : new_n2984_ = 1'b1;
default : new_n2984_ = 1'b0;
endcase
casez ({new_n166_, new_n309_, new_n767_})
3'b11? : new_n2985_ = 1'b1;
3'b??1 : new_n2985_ = 1'b1;
default : new_n2985_ = 1'b0;
endcase
casez ({new_n200_, new_n251_})
2'b00 : new_n2986_ = 1'b1;
default : new_n2986_ = 1'b0;
endcase
casez ({new_n3514_, new_n767_})
2'b1? : new_n2987_ = 1'b1;
2'b?1 : new_n2987_ = 1'b1;
default : new_n2987_ = 1'b0;
endcase
casez ({new_n196_, new_n254_})
2'b00 : new_n2988_ = 1'b1;
default : new_n2988_ = 1'b0;
endcase
casez ({new_n95_, new_n159_, new_n191_, new_n486_})
4'b11?? : new_n2989_ = 1'b1;
4'b??11 : new_n2989_ = 1'b1;
default : new_n2989_ = 1'b0;
endcase
casez ({new_n237_, new_n251_})
2'b00 : new_n2990_ = 1'b1;
default : new_n2990_ = 1'b0;
endcase
casez ({new_n182_, new_n240_, new_n201_, new_n255_})
4'b11?? : new_n2991_ = 1'b1;
4'b??11 : new_n2991_ = 1'b1;
default : new_n2991_ = 1'b0;
endcase
casez ({new_n150_, new_n488_})
2'b00 : new_n2992_ = 1'b1;
default : new_n2992_ = 1'b0;
endcase
casez ({new_n3431_, new_n222_, new_n488_})
3'b1?? : new_n2993_ = 1'b1;
3'b?11 : new_n2993_ = 1'b1;
default : new_n2993_ = 1'b0;
endcase
casez ({new_n154_, new_n284_, new_n158_, new_n488_})
4'b11?? : new_n2994_ = 1'b1;
4'b??11 : new_n2994_ = 1'b1;
default : new_n2994_ = 1'b0;
endcase
casez ({new_n169_, new_n177_, new_n170_, new_n488_})
4'b11?? : new_n2995_ = 1'b1;
4'b??11 : new_n2995_ = 1'b1;
default : new_n2995_ = 1'b0;
endcase
casez ({new_n216_, new_n247_, new_n437_, new_n488_})
4'b11?? : new_n2996_ = 1'b1;
4'b??11 : new_n2996_ = 1'b1;
default : new_n2996_ = 1'b0;
endcase
casez ({new_n145_, new_n255_})
2'b00 : new_n2997_ = 1'b1;
default : new_n2997_ = 1'b0;
endcase
casez ({u[1], new_n488_, new_n156_})
3'b01? : new_n2998_ = 1'b1;
3'b??1 : new_n2998_ = 1'b1;
default : new_n2998_ = 1'b0;
endcase
casez ({new_n3484_, new_n187_, new_n488_})
3'b1?? : new_n2999_ = 1'b1;
3'b?11 : new_n2999_ = 1'b1;
default : new_n2999_ = 1'b0;
endcase
casez ({new_n204_, new_n489_, new_n284_, new_n338_})
4'b11?? : new_n3000_ = 1'b1;
4'b??11 : new_n3000_ = 1'b1;
default : new_n3000_ = 1'b0;
endcase
casez ({new_n235_, new_n255_})
2'b00 : new_n3001_ = 1'b1;
default : new_n3001_ = 1'b0;
endcase
casez ({new_n96_, new_n135_, new_n101_, new_n143_})
4'b11?? : new_n3002_ = 1'b1;
4'b??11 : new_n3002_ = 1'b1;
default : new_n3002_ = 1'b0;
endcase
casez ({new_n142_, new_n170_, new_n3327_})
3'b11? : new_n3003_ = 1'b1;
3'b??1 : new_n3003_ = 1'b1;
default : new_n3003_ = 1'b0;
endcase
casez ({u[2], new_n85_, new_n143_})
3'b01? : new_n3004_ = 1'b1;
3'b??1 : new_n3004_ = 1'b1;
default : new_n3004_ = 1'b0;
endcase
casez ({new_n3458_, new_n237_})
2'b1? : new_n3005_ = 1'b1;
2'b?1 : new_n3005_ = 1'b1;
default : new_n3005_ = 1'b0;
endcase
casez ({new_n86_, new_n258_})
2'b00 : new_n3006_ = 1'b1;
default : new_n3006_ = 1'b0;
endcase
casez ({new_n204_, new_n258_})
2'b00 : new_n3007_ = 1'b1;
default : new_n3007_ = 1'b0;
endcase
casez ({new_n3330_, new_n187_, new_n198_})
3'b1?? : new_n3008_ = 1'b1;
3'b?11 : new_n3008_ = 1'b1;
default : new_n3008_ = 1'b0;
endcase
casez ({new_n140_, new_n144_})
2'b00 : new_n3009_ = 1'b1;
default : new_n3009_ = 1'b0;
endcase
casez ({new_n189_, new_n500_})
2'b00 : new_n3010_ = 1'b1;
default : new_n3010_ = 1'b0;
endcase
casez ({new_n158_, new_n214_, new_n3459_})
3'b11? : new_n3011_ = 1'b1;
3'b??1 : new_n3011_ = 1'b1;
default : new_n3011_ = 1'b0;
endcase
casez ({new_n3598_, new_n3460_})
2'b1? : new_n3012_ = 1'b1;
2'b?1 : new_n3012_ = 1'b1;
default : new_n3012_ = 1'b0;
endcase
casez ({new_n3527_, new_n210_, new_n261_})
3'b1?? : new_n3013_ = 1'b1;
3'b?11 : new_n3013_ = 1'b1;
default : new_n3013_ = 1'b0;
endcase
casez ({new_n222_, new_n262_})
2'b00 : new_n3014_ = 1'b1;
default : new_n3014_ = 1'b0;
endcase
casez ({new_n151_, new_n190_, new_n191_, new_n262_})
4'b11?? : new_n3015_ = 1'b1;
4'b??11 : new_n3015_ = 1'b1;
default : new_n3015_ = 1'b0;
endcase
casez ({new_n219_, new_n262_, new_n244_, new_n249_})
4'b11?? : new_n3016_ = 1'b1;
4'b??11 : new_n3016_ = 1'b1;
default : new_n3016_ = 1'b0;
endcase
casez ({new_n173_, new_n262_})
2'b00 : new_n3017_ = 1'b1;
default : new_n3017_ = 1'b0;
endcase
casez ({new_n144_, new_n508_, new_n3349_})
3'b11? : new_n3018_ = 1'b1;
3'b??1 : new_n3018_ = 1'b1;
default : new_n3018_ = 1'b0;
endcase
casez ({new_n167_, new_n356_, new_n192_, new_n508_})
4'b11?? : new_n3019_ = 1'b1;
4'b??11 : new_n3019_ = 1'b1;
default : new_n3019_ = 1'b0;
endcase
casez ({new_n115_, new_n148_})
2'b00 : new_n3020_ = 1'b1;
default : new_n3020_ = 1'b0;
endcase
casez ({new_n187_, new_n264_, new_n200_, new_n209_})
4'b11?? : new_n3021_ = 1'b1;
4'b??11 : new_n3021_ = 1'b1;
default : new_n3021_ = 1'b0;
endcase
casez ({new_n3571_, new_n86_, new_n509_})
3'b1?? : new_n3022_ = 1'b1;
3'b?11 : new_n3022_ = 1'b1;
default : new_n3022_ = 1'b0;
endcase
casez ({new_n3513_, new_n3340_})
2'b1? : new_n3023_ = 1'b1;
2'b?1 : new_n3023_ = 1'b1;
default : new_n3023_ = 1'b0;
endcase
casez ({new_n3376_, new_n166_, new_n509_})
3'b1?? : new_n3024_ = 1'b1;
3'b?11 : new_n3024_ = 1'b1;
default : new_n3024_ = 1'b0;
endcase
casez ({new_n150_, new_n264_})
2'b00 : new_n3025_ = 1'b1;
default : new_n3025_ = 1'b0;
endcase
casez ({new_n85_, new_n97_, new_n148_})
3'b11? : new_n3026_ = 1'b1;
3'b??1 : new_n3026_ = 1'b1;
default : new_n3026_ = 1'b0;
endcase
casez ({new_n88_, new_n150_, new_n223_, new_n264_})
4'b11?? : new_n3027_ = 1'b1;
4'b??11 : new_n3027_ = 1'b1;
default : new_n3027_ = 1'b0;
endcase
casez ({new_n139_, new_n148_})
2'b00 : new_n3028_ = 1'b1;
default : new_n3028_ = 1'b0;
endcase
casez ({new_n173_, new_n230_, new_n258_, new_n266_})
4'b11?? : new_n3029_ = 1'b1;
4'b??11 : new_n3029_ = 1'b1;
default : new_n3029_ = 1'b0;
endcase
casez ({new_n205_, new_n266_})
2'b00 : new_n3030_ = 1'b1;
default : new_n3030_ = 1'b0;
endcase
casez ({v[0], new_n150_, new_n100_, new_n139_})
4'b11?? : new_n3031_ = 1'b1;
4'b??11 : new_n3031_ = 1'b1;
default : new_n3031_ = 1'b0;
endcase
casez ({new_n217_, new_n266_})
2'b00 : new_n3032_ = 1'b1;
default : new_n3032_ = 1'b0;
endcase
casez ({new_n145_, new_n176_, new_n204_, new_n266_})
4'b11?? : new_n3033_ = 1'b1;
4'b??11 : new_n3033_ = 1'b1;
default : new_n3033_ = 1'b0;
endcase
casez ({new_n244_, new_n266_})
2'b00 : new_n3034_ = 1'b1;
default : new_n3034_ = 1'b0;
endcase
casez ({new_n80_, new_n190_, new_n216_, new_n266_})
4'b11?? : new_n3035_ = 1'b1;
4'b??11 : new_n3035_ = 1'b1;
default : new_n3035_ = 1'b0;
endcase
casez ({new_n145_, new_n201_, new_n151_, new_n522_})
4'b11?? : new_n3036_ = 1'b1;
4'b??11 : new_n3036_ = 1'b1;
default : new_n3036_ = 1'b0;
endcase
casez ({new_n94_, new_n182_, new_n215_, new_n522_})
4'b11?? : new_n3037_ = 1'b1;
4'b??11 : new_n3037_ = 1'b1;
default : new_n3037_ = 1'b0;
endcase
casez ({x[2], new_n153_, new_n86_, new_n98_})
4'b01?? : new_n3038_ = 1'b1;
4'b??11 : new_n3038_ = 1'b1;
default : new_n3038_ = 1'b0;
endcase
casez ({x[1], new_n98_, new_n153_})
3'b01? : new_n3039_ = 1'b1;
3'b??1 : new_n3039_ = 1'b1;
default : new_n3039_ = 1'b0;
endcase
casez ({new_n3609_, new_n3465_})
2'b1? : new_n3040_ = 1'b1;
2'b?1 : new_n3040_ = 1'b1;
default : new_n3040_ = 1'b0;
endcase
casez ({new_n104_, new_n153_, new_n133_})
3'b11? : new_n3041_ = 1'b1;
3'b??1 : new_n3041_ = 1'b1;
default : new_n3041_ = 1'b0;
endcase
casez ({new_n80_, new_n261_, new_n363_, new_n530_})
4'b11?? : new_n3042_ = 1'b1;
4'b??11 : new_n3042_ = 1'b1;
default : new_n3042_ = 1'b0;
endcase
casez ({new_n88_, new_n530_, new_n167_, new_n522_})
4'b11?? : new_n3043_ = 1'b1;
4'b??11 : new_n3043_ = 1'b1;
default : new_n3043_ = 1'b0;
endcase
casez ({x[2], new_n273_, v[1], new_n152_})
4'b01?? : new_n3044_ = 1'b1;
4'b??11 : new_n3044_ = 1'b1;
default : new_n3044_ = 1'b0;
endcase
casez ({new_n161_, new_n273_, new_n3517_})
3'b11? : new_n3045_ = 1'b1;
3'b??1 : new_n3045_ = 1'b1;
default : new_n3045_ = 1'b0;
endcase
casez ({new_n3467_, new_n3567_})
2'b1? : new_n3046_ = 1'b1;
2'b?1 : new_n3046_ = 1'b1;
default : new_n3046_ = 1'b0;
endcase
casez ({new_n97_, new_n177_, new_n204_, new_n274_})
4'b11?? : new_n3047_ = 1'b1;
4'b??11 : new_n3047_ = 1'b1;
default : new_n3047_ = 1'b0;
endcase
casez ({new_n209_, new_n274_})
2'b00 : new_n3048_ = 1'b1;
default : new_n3048_ = 1'b0;
endcase
casez ({new_n162_, new_n274_})
2'b00 : new_n3049_ = 1'b1;
default : new_n3049_ = 1'b0;
endcase
casez ({new_n104_, new_n214_, new_n3350_})
3'b11? : new_n3050_ = 1'b1;
3'b??1 : new_n3050_ = 1'b1;
default : new_n3050_ = 1'b0;
endcase
casez ({new_n207_, new_n274_})
2'b00 : new_n3051_ = 1'b1;
default : new_n3051_ = 1'b0;
endcase
casez ({new_n148_, new_n210_, new_n3352_})
3'b11? : new_n3052_ = 1'b1;
3'b??1 : new_n3052_ = 1'b1;
default : new_n3052_ = 1'b0;
endcase
casez ({x[2], new_n162_, new_n275_})
3'b11? : new_n3053_ = 1'b1;
3'b??1 : new_n3053_ = 1'b1;
default : new_n3053_ = 1'b0;
endcase
casez ({new_n155_, new_n821_})
2'b00 : new_n3054_ = 1'b1;
default : new_n3054_ = 1'b0;
endcase
casez ({new_n142_, new_n247_, new_n154_, new_n822_})
4'b11?? : new_n3055_ = 1'b1;
4'b??11 : new_n3055_ = 1'b1;
default : new_n3055_ = 1'b0;
endcase
casez ({new_n3449_, new_n488_, new_n822_})
3'b1?? : new_n3056_ = 1'b1;
3'b?11 : new_n3056_ = 1'b1;
default : new_n3056_ = 1'b0;
endcase
casez ({new_n3607_, new_n264_, new_n278_})
3'b1?? : new_n3057_ = 1'b1;
3'b?11 : new_n3057_ = 1'b1;
default : new_n3057_ = 1'b0;
endcase
casez ({new_n144_, new_n278_, new_n161_, new_n221_})
4'b11?? : new_n3058_ = 1'b1;
4'b??11 : new_n3058_ = 1'b1;
default : new_n3058_ = 1'b0;
endcase
casez ({new_n207_, new_n279_, new_n216_, new_n235_})
4'b11?? : new_n3059_ = 1'b1;
4'b??11 : new_n3059_ = 1'b1;
default : new_n3059_ = 1'b0;
endcase
casez ({new_n3532_, new_n251_, new_n279_})
3'b1?? : new_n3060_ = 1'b1;
3'b?11 : new_n3060_ = 1'b1;
default : new_n3060_ = 1'b0;
endcase
casez ({new_n160_, new_n261_, new_n187_, new_n279_})
4'b11?? : new_n3061_ = 1'b1;
4'b??11 : new_n3061_ = 1'b1;
default : new_n3061_ = 1'b0;
endcase
casez ({new_n89_, new_n160_})
2'b00 : new_n3062_ = 1'b1;
default : new_n3062_ = 1'b0;
endcase
casez ({new_n173_, new_n258_, new_n192_, new_n279_})
4'b11?? : new_n3063_ = 1'b1;
4'b??11 : new_n3063_ = 1'b1;
default : new_n3063_ = 1'b0;
endcase
casez ({new_n222_, new_n279_})
2'b00 : new_n3064_ = 1'b1;
default : new_n3064_ = 1'b0;
endcase
casez ({new_n3473_, new_n123_, new_n254_})
3'b1?? : new_n3065_ = 1'b1;
3'b?11 : new_n3065_ = 1'b1;
default : new_n3065_ = 1'b0;
endcase
casez ({new_n79_, new_n160_, new_n3342_})
3'b11? : new_n3066_ = 1'b1;
3'b??1 : new_n3066_ = 1'b1;
default : new_n3066_ = 1'b0;
endcase
casez ({new_n167_, new_n281_})
2'b00 : new_n3067_ = 1'b1;
default : new_n3067_ = 1'b0;
endcase
casez ({new_n148_, new_n281_, new_n3488_})
3'b11? : new_n3068_ = 1'b1;
3'b??1 : new_n3068_ = 1'b1;
default : new_n3068_ = 1'b0;
endcase
casez ({new_n88_, new_n161_})
2'b00 : new_n3069_ = 1'b1;
default : new_n3069_ = 1'b0;
endcase
casez ({new_n142_, new_n281_, new_n169_, new_n192_})
4'b11?? : new_n3070_ = 1'b1;
4'b??11 : new_n3070_ = 1'b1;
default : new_n3070_ = 1'b0;
endcase
casez ({new_n3608_, new_n3355_})
2'b1? : new_n3071_ = 1'b1;
2'b?1 : new_n3071_ = 1'b1;
default : new_n3071_ = 1'b0;
endcase
casez ({new_n90_, new_n158_, new_n191_, new_n549_})
4'b11?? : new_n3072_ = 1'b1;
4'b??11 : new_n3072_ = 1'b1;
default : new_n3072_ = 1'b0;
endcase
casez ({new_n82_, new_n91_, new_n285_})
3'b10? : new_n3073_ = 1'b1;
3'b??1 : new_n3073_ = 1'b1;
default : new_n3073_ = 1'b0;
endcase
casez ({new_n228_, new_n285_})
2'b00 : new_n3074_ = 1'b1;
default : new_n3074_ = 1'b0;
endcase
casez ({new_n166_, new_n279_, new_n204_, new_n285_})
4'b11?? : new_n3075_ = 1'b1;
4'b??11 : new_n3075_ = 1'b1;
default : new_n3075_ = 1'b0;
endcase
casez ({new_n173_, new_n184_, new_n199_, new_n285_})
4'b11?? : new_n3076_ = 1'b1;
4'b??11 : new_n3076_ = 1'b1;
default : new_n3076_ = 1'b0;
endcase
casez ({new_n80_, new_n173_, new_n3356_})
3'b11? : new_n3077_ = 1'b1;
3'b??1 : new_n3077_ = 1'b1;
default : new_n3077_ = 1'b0;
endcase
casez ({new_n196_, new_n363_, new_n199_, new_n1257_})
4'b11?? : new_n3078_ = 1'b1;
4'b??11 : new_n3078_ = 1'b1;
default : new_n3078_ = 1'b0;
endcase
casez ({new_n107_, new_n1258_, new_n242_})
3'b01? : new_n3079_ = 1'b1;
3'b??1 : new_n3079_ = 1'b1;
default : new_n3079_ = 1'b0;
endcase
casez ({new_n169_, new_n201_, new_n243_, new_n1258_})
4'b11?? : new_n3080_ = 1'b1;
4'b??11 : new_n3080_ = 1'b1;
default : new_n3080_ = 1'b0;
endcase
casez ({new_n3446_, new_n321_, new_n1262_})
3'b1?? : new_n3081_ = 1'b1;
3'b?10 : new_n3081_ = 1'b1;
default : new_n3081_ = 1'b0;
endcase
casez ({new_n93_, new_n1262_, new_n293_})
3'b10? : new_n3082_ = 1'b1;
3'b??1 : new_n3082_ = 1'b1;
default : new_n3082_ = 1'b0;
endcase
casez ({new_n139_, new_n237_, new_n1266_})
3'b11? : new_n3083_ = 1'b1;
3'b??1 : new_n3083_ = 1'b1;
default : new_n3083_ = 1'b0;
endcase
casez ({new_n167_, new_n1267_})
2'b00 : new_n3084_ = 1'b1;
default : new_n3084_ = 1'b0;
endcase
casez ({new_n89_, new_n116_, new_n3585_})
3'b01? : new_n3085_ = 1'b1;
3'b??1 : new_n3085_ = 1'b1;
default : new_n3085_ = 1'b0;
endcase
casez ({new_n3572_, new_n565_})
2'b1? : new_n3086_ = 1'b1;
2'b?1 : new_n3086_ = 1'b1;
default : new_n3086_ = 1'b0;
endcase
casez ({new_n3440_, new_n565_})
2'b1? : new_n3087_ = 1'b1;
2'b?1 : new_n3087_ = 1'b1;
default : new_n3087_ = 1'b0;
endcase
casez ({new_n158_, new_n167_})
2'b00 : new_n3088_ = 1'b1;
default : new_n3088_ = 1'b0;
endcase
casez ({x[1], new_n293_, new_n101_, new_n163_})
4'b01?? : new_n3089_ = 1'b1;
4'b??11 : new_n3089_ = 1'b1;
default : new_n3089_ = 1'b0;
endcase
casez ({new_n80_, new_n251_, new_n93_, new_n293_})
4'b11?? : new_n3090_ = 1'b1;
4'b??11 : new_n3090_ = 1'b1;
default : new_n3090_ = 1'b0;
endcase
casez ({new_n3322_, new_n3363_})
2'b1? : new_n3091_ = 1'b1;
2'b?1 : new_n3091_ = 1'b1;
default : new_n3091_ = 1'b0;
endcase
casez ({new_n235_, new_n299_})
2'b00 : new_n3092_ = 1'b1;
default : new_n3092_ = 1'b0;
endcase
casez ({new_n142_, new_n255_, new_n153_, new_n299_})
4'b11?? : new_n3093_ = 1'b1;
4'b??11 : new_n3093_ = 1'b1;
default : new_n3093_ = 1'b0;
endcase
casez ({new_n142_, new_n221_, new_n214_, new_n299_})
4'b11?? : new_n3094_ = 1'b1;
4'b??11 : new_n3094_ = 1'b1;
default : new_n3094_ = 1'b0;
endcase
casez ({new_n3563_, new_n129_, new_n170_})
3'b1?? : new_n3095_ = 1'b1;
3'b?11 : new_n3095_ = 1'b1;
default : new_n3095_ = 1'b0;
endcase
casez ({new_n89_, new_n299_, new_n173_})
3'b01? : new_n3096_ = 1'b1;
3'b??1 : new_n3096_ = 1'b1;
default : new_n3096_ = 1'b0;
endcase
casez ({new_n144_, new_n300_, new_n182_, new_n222_})
4'b11?? : new_n3097_ = 1'b1;
4'b??11 : new_n3097_ = 1'b1;
default : new_n3097_ = 1'b0;
endcase
casez ({new_n215_, new_n300_})
2'b00 : new_n3098_ = 1'b1;
default : new_n3098_ = 1'b0;
endcase
casez ({new_n145_, new_n173_})
2'b00 : new_n3099_ = 1'b1;
default : new_n3099_ = 1'b0;
endcase
casez ({new_n3474_, new_n3367_})
2'b1? : new_n3100_ = 1'b1;
2'b?1 : new_n3100_ = 1'b1;
default : new_n3100_ = 1'b0;
endcase
casez ({new_n254_, new_n305_})
2'b00 : new_n3101_ = 1'b1;
default : new_n3101_ = 1'b0;
endcase
casez ({new_n3352_, new_n169_, new_n305_})
3'b1?? : new_n3102_ = 1'b1;
3'b?11 : new_n3102_ = 1'b1;
default : new_n3102_ = 1'b0;
endcase
casez ({u[2], new_n161_, new_n176_})
3'b11? : new_n3103_ = 1'b1;
3'b??1 : new_n3103_ = 1'b1;
default : new_n3103_ = 1'b0;
endcase
casez ({new_n207_, new_n309_})
2'b00 : new_n3104_ = 1'b1;
default : new_n3104_ = 1'b0;
endcase
casez ({new_n3522_, new_n86_, new_n309_})
3'b1?? : new_n3105_ = 1'b1;
3'b?11 : new_n3105_ = 1'b1;
default : new_n3105_ = 1'b0;
endcase
casez ({new_n215_, new_n597_, new_n247_, new_n305_})
4'b11?? : new_n3106_ = 1'b1;
4'b??11 : new_n3106_ = 1'b1;
default : new_n3106_ = 1'b0;
endcase
casez ({new_n170_, new_n309_, new_n3388_})
3'b11? : new_n3107_ = 1'b1;
3'b??1 : new_n3107_ = 1'b1;
default : new_n3107_ = 1'b0;
endcase
casez ({new_n3498_, new_n237_, new_n598_})
3'b1?? : new_n3108_ = 1'b1;
3'b?11 : new_n3108_ = 1'b1;
default : new_n3108_ = 1'b0;
endcase
casez ({y[2], new_n255_, new_n83_, new_n598_})
4'b11?? : new_n3109_ = 1'b1;
4'b??11 : new_n3109_ = 1'b1;
default : new_n3109_ = 1'b0;
endcase
casez ({new_n178_, new_n598_, new_n229_, new_n522_})
4'b11?? : new_n3110_ = 1'b1;
4'b??11 : new_n3110_ = 1'b1;
default : new_n3110_ = 1'b0;
endcase
casez ({new_n142_, new_n215_, new_n143_, new_n599_})
4'b11?? : new_n3111_ = 1'b1;
4'b??11 : new_n3111_ = 1'b1;
default : new_n3111_ = 1'b0;
endcase
casez ({new_n158_, new_n178_})
2'b00 : new_n3112_ = 1'b1;
default : new_n3112_ = 1'b0;
endcase
casez ({new_n213_, new_n313_})
2'b00 : new_n3113_ = 1'b1;
default : new_n3113_ = 1'b0;
endcase
casez ({new_n170_, new_n218_, new_n204_, new_n313_})
4'b11?? : new_n3114_ = 1'b1;
4'b??11 : new_n3114_ = 1'b1;
default : new_n3114_ = 1'b0;
endcase
casez ({new_n3421_, new_n3373_})
2'b1? : new_n3115_ = 1'b1;
2'b?1 : new_n3115_ = 1'b1;
default : new_n3115_ = 1'b0;
endcase
casez ({new_n161_, new_n275_, new_n3374_})
3'b11? : new_n3116_ = 1'b1;
3'b??1 : new_n3116_ = 1'b1;
default : new_n3116_ = 1'b0;
endcase
casez ({new_n3375_, new_n150_})
2'b1? : new_n3117_ = 1'b1;
2'b?1 : new_n3117_ = 1'b1;
default : new_n3117_ = 1'b0;
endcase
casez ({new_n148_, new_n170_, new_n158_, new_n317_})
4'b11?? : new_n3118_ = 1'b1;
4'b??11 : new_n3118_ = 1'b1;
default : new_n3118_ = 1'b0;
endcase
casez ({new_n249_, new_n316_})
2'b00 : new_n3119_ = 1'b1;
default : new_n3119_ = 1'b0;
endcase
casez ({new_n3377_, new_n209_, new_n254_})
3'b1?? : new_n3120_ = 1'b1;
3'b?11 : new_n3120_ = 1'b1;
default : new_n3120_ = 1'b0;
endcase
casez ({new_n115_, new_n317_})
2'b00 : new_n3121_ = 1'b1;
default : new_n3121_ = 1'b0;
endcase
casez ({new_n204_, new_n317_, new_n248_, new_n309_})
4'b11?? : new_n3122_ = 1'b1;
4'b??11 : new_n3122_ = 1'b1;
default : new_n3122_ = 1'b0;
endcase
casez ({new_n98_, new_n2495_, new_n1799_})
3'b11? : new_n3123_ = 1'b1;
3'b??1 : new_n3123_ = 1'b1;
default : new_n3123_ = 1'b0;
endcase
casez ({new_n166_, new_n209_, new_n167_, new_n317_})
4'b11?? : new_n3124_ = 1'b1;
4'b??11 : new_n3124_ = 1'b1;
default : new_n3124_ = 1'b0;
endcase
casez ({new_n109_, new_n2497_, new_n230_})
3'b01? : new_n3125_ = 1'b1;
3'b??1 : new_n3125_ = 1'b1;
default : new_n3125_ = 1'b0;
endcase
casez ({new_n82_, new_n150_, new_n155_, new_n2500_})
4'b11?? : new_n3126_ = 1'b1;
4'b??10 : new_n3126_ = 1'b1;
default : new_n3126_ = 1'b0;
endcase
casez ({new_n199_, new_n2502_})
2'b00 : new_n3127_ = 1'b1;
default : new_n3127_ = 1'b0;
endcase
casez ({new_n167_, new_n241_, new_n242_, new_n317_})
4'b11?? : new_n3128_ = 1'b1;
4'b??11 : new_n3128_ = 1'b1;
default : new_n3128_ = 1'b0;
endcase
casez ({new_n158_, new_n182_})
2'b00 : new_n3129_ = 1'b1;
default : new_n3129_ = 1'b0;
endcase
casez ({new_n1542_, new_n2507_})
2'b00 : new_n3130_ = 1'b1;
default : new_n3130_ = 1'b0;
endcase
casez ({new_n238_, new_n2508_})
2'b00 : new_n3131_ = 1'b1;
default : new_n3131_ = 1'b0;
endcase
casez ({new_n307_, new_n2510_})
2'b00 : new_n3132_ = 1'b1;
default : new_n3132_ = 1'b0;
endcase
casez ({new_n98_, new_n255_, new_n2512_})
3'b01? : new_n3133_ = 1'b1;
3'b??1 : new_n3133_ = 1'b1;
default : new_n3133_ = 1'b0;
endcase
casez ({new_n189_, new_n250_, new_n194_, new_n2513_})
4'b11?? : new_n3134_ = 1'b1;
4'b??11 : new_n3134_ = 1'b1;
default : new_n3134_ = 1'b0;
endcase
casez ({new_n81_, new_n2514_})
2'b00 : new_n3135_ = 1'b1;
default : new_n3135_ = 1'b0;
endcase
casez ({new_n94_, new_n210_, new_n217_, new_n2515_})
4'b11?? : new_n3136_ = 1'b1;
4'b??11 : new_n3136_ = 1'b1;
default : new_n3136_ = 1'b0;
endcase
casez ({new_n169_, new_n318_, new_n205_, new_n216_})
4'b11?? : new_n3137_ = 1'b1;
4'b??11 : new_n3137_ = 1'b1;
default : new_n3137_ = 1'b0;
endcase
casez ({new_n123_, new_n2518_})
2'b00 : new_n3138_ = 1'b1;
default : new_n3138_ = 1'b0;
endcase
casez ({new_n199_, new_n2519_})
2'b00 : new_n3139_ = 1'b1;
default : new_n3139_ = 1'b0;
endcase
casez ({u[2], new_n159_, new_n2521_})
3'b11? : new_n3140_ = 1'b1;
3'b??1 : new_n3140_ = 1'b1;
default : new_n3140_ = 1'b0;
endcase
casez ({new_n178_, new_n183_})
2'b00 : new_n3141_ = 1'b1;
default : new_n3141_ = 1'b0;
endcase
casez ({new_n216_, new_n299_, new_n244_, new_n321_})
4'b11?? : new_n3142_ = 1'b1;
4'b??11 : new_n3142_ = 1'b1;
default : new_n3142_ = 1'b0;
endcase
casez ({new_n139_, new_n321_})
2'b00 : new_n3143_ = 1'b1;
default : new_n3143_ = 1'b0;
endcase
casez ({new_n142_, new_n210_, new_n3379_})
3'b11? : new_n3144_ = 1'b1;
3'b??1 : new_n3144_ = 1'b1;
default : new_n3144_ = 1'b0;
endcase
casez ({y[1], new_n118_, new_n3380_})
3'b01? : new_n3145_ = 1'b1;
3'b??1 : new_n3145_ = 1'b1;
default : new_n3145_ = 1'b0;
endcase
casez ({new_n3429_, new_n261_, new_n321_})
3'b1?? : new_n3146_ = 1'b1;
3'b?11 : new_n3146_ = 1'b1;
default : new_n3146_ = 1'b0;
endcase
casez ({new_n182_, new_n184_})
2'b00 : new_n3147_ = 1'b1;
default : new_n3147_ = 1'b0;
endcase
casez ({new_n177_, new_n184_})
2'b00 : new_n3148_ = 1'b1;
default : new_n3148_ = 1'b0;
endcase
casez ({new_n3361_, new_n93_, new_n184_})
3'b1?? : new_n3149_ = 1'b1;
3'b?11 : new_n3149_ = 1'b1;
default : new_n3149_ = 1'b0;
endcase
casez ({new_n196_, new_n260_, new_n204_, new_n923_})
4'b11?? : new_n3150_ = 1'b1;
4'b??11 : new_n3150_ = 1'b1;
default : new_n3150_ = 1'b0;
endcase
casez ({new_n3333_, new_n237_, new_n923_})
3'b1?? : new_n3151_ = 1'b1;
3'b?11 : new_n3151_ = 1'b1;
default : new_n3151_ = 1'b0;
endcase
casez ({new_n299_, new_n924_})
2'b00 : new_n3152_ = 1'b1;
default : new_n3152_ = 1'b0;
endcase
casez ({new_n96_, new_n118_, new_n248_, new_n328_})
4'b11?? : new_n3153_ = 1'b1;
4'b??11 : new_n3153_ = 1'b1;
default : new_n3153_ = 1'b0;
endcase
casez ({new_n145_, new_n328_, new_n217_, new_n287_})
4'b11?? : new_n3154_ = 1'b1;
4'b??11 : new_n3154_ = 1'b1;
default : new_n3154_ = 1'b0;
endcase
casez ({new_n293_, new_n926_})
2'b00 : new_n3155_ = 1'b1;
default : new_n3155_ = 1'b0;
endcase
casez ({new_n3501_, new_n131_, new_n184_})
3'b1?? : new_n3156_ = 1'b1;
3'b?11 : new_n3156_ = 1'b1;
default : new_n3156_ = 1'b0;
endcase
casez ({new_n173_, new_n332_, new_n3359_})
3'b11? : new_n3157_ = 1'b1;
3'b??1 : new_n3157_ = 1'b1;
default : new_n3157_ = 1'b0;
endcase
casez ({new_n129_, new_n332_, new_n241_, new_n262_})
4'b11?? : new_n3158_ = 1'b1;
4'b??11 : new_n3158_ = 1'b1;
default : new_n3158_ = 1'b0;
endcase
casez ({new_n169_, new_n332_})
2'b00 : new_n3159_ = 1'b1;
default : new_n3159_ = 1'b0;
endcase
casez ({new_n95_, new_n211_, new_n137_, new_n332_})
4'b11?? : new_n3160_ = 1'b1;
4'b??11 : new_n3160_ = 1'b1;
default : new_n3160_ = 1'b0;
endcase
casez ({new_n129_, new_n189_})
2'b00 : new_n3161_ = 1'b1;
default : new_n3161_ = 1'b0;
endcase
casez ({u[0], new_n231_, new_n88_, new_n337_})
4'b01?? : new_n3162_ = 1'b1;
4'b??01 : new_n3162_ = 1'b1;
default : new_n3162_ = 1'b0;
endcase
casez ({new_n100_, new_n153_, new_n338_})
3'b11? : new_n3163_ = 1'b1;
3'b??1 : new_n3163_ = 1'b1;
default : new_n3163_ = 1'b0;
endcase
casez ({new_n118_, new_n194_})
2'b00 : new_n3164_ = 1'b1;
default : new_n3164_ = 1'b0;
endcase
casez ({new_n3508_, new_n118_, new_n173_})
3'b1?? : new_n3165_ = 1'b1;
3'b?11 : new_n3165_ = 1'b1;
default : new_n3165_ = 1'b0;
endcase
casez ({new_n160_, new_n309_, new_n177_, new_n343_})
4'b11?? : new_n3166_ = 1'b1;
4'b??11 : new_n3166_ = 1'b1;
default : new_n3166_ = 1'b0;
endcase
casez ({new_n3485_, new_n3390_})
2'b1? : new_n3167_ = 1'b1;
2'b?1 : new_n3167_ = 1'b1;
default : new_n3167_ = 1'b0;
endcase
casez ({new_n3589_, new_n99_, new_n343_})
3'b1?? : new_n3168_ = 1'b1;
3'b?01 : new_n3168_ = 1'b1;
default : new_n3168_ = 1'b0;
endcase
casez ({new_n3390_, new_n3457_})
2'b1? : new_n3169_ = 1'b1;
2'b?1 : new_n3169_ = 1'b1;
default : new_n3169_ = 1'b0;
endcase
casez ({new_n176_, new_n343_, new_n194_, new_n224_})
4'b11?? : new_n3170_ = 1'b1;
4'b??11 : new_n3170_ = 1'b1;
default : new_n3170_ = 1'b0;
endcase
casez ({new_n85_, new_n196_})
2'b00 : new_n3171_ = 1'b1;
default : new_n3171_ = 1'b0;
endcase
casez ({new_n208_, new_n264_, new_n211_, new_n344_})
4'b11?? : new_n3172_ = 1'b1;
4'b??11 : new_n3172_ = 1'b1;
default : new_n3172_ = 1'b0;
endcase
casez ({new_n161_, new_n344_})
2'b00 : new_n3173_ = 1'b1;
default : new_n3173_ = 1'b0;
endcase
casez ({new_n3392_, new_n204_, new_n217_})
3'b1?? : new_n3174_ = 1'b1;
3'b?11 : new_n3174_ = 1'b1;
default : new_n3174_ = 1'b0;
endcase
casez ({new_n89_, new_n150_, new_n3395_})
3'b11? : new_n3175_ = 1'b1;
3'b??1 : new_n3175_ = 1'b1;
default : new_n3175_ = 1'b0;
endcase
casez ({v[2], new_n115_, new_n3510_})
3'b01? : new_n3176_ = 1'b1;
3'b??1 : new_n3176_ = 1'b1;
default : new_n3176_ = 1'b0;
endcase
casez ({new_n191_, new_n199_})
2'b00 : new_n3177_ = 1'b1;
default : new_n3177_ = 1'b0;
endcase
casez ({new_n158_, new_n200_})
2'b00 : new_n3178_ = 1'b1;
default : new_n3178_ = 1'b0;
endcase
casez ({new_n3515_, new_n347_})
2'b1? : new_n3179_ = 1'b1;
2'b?1 : new_n3179_ = 1'b1;
default : new_n3179_ = 1'b0;
endcase
casez ({x[1], new_n237_, u[2], new_n347_})
4'b11?? : new_n3180_ = 1'b1;
4'b??01 : new_n3180_ = 1'b1;
default : new_n3180_ = 1'b0;
endcase
casez ({new_n3368_, new_n241_, new_n347_})
3'b1?? : new_n3181_ = 1'b1;
3'b?11 : new_n3181_ = 1'b1;
default : new_n3181_ = 1'b0;
endcase
casez ({x[1], new_n301_, new_n347_})
3'b01? : new_n3182_ = 1'b1;
3'b??1 : new_n3182_ = 1'b1;
default : new_n3182_ = 1'b0;
endcase
casez ({new_n3399_, new_n148_, new_n184_})
3'b1?? : new_n3183_ = 1'b1;
3'b?11 : new_n3183_ = 1'b1;
default : new_n3183_ = 1'b0;
endcase
casez ({new_n104_, new_n356_, new_n3369_})
3'b11? : new_n3184_ = 1'b1;
3'b??1 : new_n3184_ = 1'b1;
default : new_n3184_ = 1'b0;
endcase
casez ({new_n150_, new_n224_, new_n3402_})
3'b11? : new_n3185_ = 1'b1;
3'b??1 : new_n3185_ = 1'b1;
default : new_n3185_ = 1'b0;
endcase
casez ({new_n153_, new_n170_, new_n158_, new_n356_})
4'b11?? : new_n3186_ = 1'b1;
4'b??11 : new_n3186_ = 1'b1;
default : new_n3186_ = 1'b0;
endcase
casez ({new_n356_, new_n358_})
2'b00 : new_n3187_ = 1'b1;
default : new_n3187_ = 1'b0;
endcase
casez ({new_n150_, new_n266_, new_n306_, new_n363_})
4'b11?? : new_n3188_ = 1'b1;
4'b??11 : new_n3188_ = 1'b1;
default : new_n3188_ = 1'b0;
endcase
casez ({x[2], new_n363_, v[1], new_n163_})
4'b11?? : new_n3189_ = 1'b1;
4'b??11 : new_n3189_ = 1'b1;
default : new_n3189_ = 1'b0;
endcase
casez ({new_n167_, new_n363_, new_n199_, new_n273_})
4'b11?? : new_n3190_ = 1'b1;
4'b??11 : new_n3190_ = 1'b1;
default : new_n3190_ = 1'b0;
endcase
casez ({new_n142_, new_n363_})
2'b00 : new_n3191_ = 1'b1;
default : new_n3191_ = 1'b0;
endcase
casez ({x[0], new_n205_, new_n3568_})
3'b01? : new_n3192_ = 1'b1;
3'b??1 : new_n3192_ = 1'b1;
default : new_n3192_ = 1'b0;
endcase
casez ({new_n3400_, new_n210_, new_n363_})
3'b1?? : new_n3193_ = 1'b1;
3'b?11 : new_n3193_ = 1'b1;
default : new_n3193_ = 1'b0;
endcase
casez ({new_n3432_, new_n3411_})
2'b1? : new_n3194_ = 1'b1;
2'b?1 : new_n3194_ = 1'b1;
default : new_n3194_ = 1'b0;
endcase
casez ({new_n3436_, new_n216_, new_n1544_})
3'b1?? : new_n3195_ = 1'b1;
3'b?11 : new_n3195_ = 1'b1;
default : new_n3195_ = 1'b0;
endcase
casez ({new_n79_, new_n151_, new_n89_, new_n1546_})
4'b11?? : new_n3196_ = 1'b1;
4'b??01 : new_n3196_ = 1'b1;
default : new_n3196_ = 1'b0;
endcase
casez ({new_n115_, new_n207_})
2'b00 : new_n3197_ = 1'b1;
default : new_n3197_ = 1'b0;
endcase
casez ({new_n3415_, new_n237_, new_n369_})
3'b1?? : new_n3198_ = 1'b1;
3'b?11 : new_n3198_ = 1'b1;
default : new_n3198_ = 1'b0;
endcase
casez ({new_n98_, new_n2915_, new_n154_})
3'b11? : new_n3199_ = 1'b1;
3'b??1 : new_n3199_ = 1'b1;
default : new_n3199_ = 1'b0;
endcase
casez ({new_n2915_, new_n2918_})
2'b01 : new_n3200_ = 1'b1;
default : new_n3200_ = 1'b0;
endcase
casez ({new_n3605_, new_n284_, new_n369_})
3'b1?? : new_n3201_ = 1'b1;
3'b?11 : new_n3201_ = 1'b1;
default : new_n3201_ = 1'b0;
endcase
casez ({new_n123_, new_n2938_})
2'b00 : new_n3202_ = 1'b1;
default : new_n3202_ = 1'b0;
endcase
casez ({new_n182_, new_n2943_})
2'b00 : new_n3203_ = 1'b1;
default : new_n3203_ = 1'b0;
endcase
casez ({new_n3328_, new_n3417_})
2'b1? : new_n3204_ = 1'b1;
2'b?1 : new_n3204_ = 1'b1;
default : new_n3204_ = 1'b0;
endcase
casez ({new_n160_, new_n2948_})
2'b00 : new_n3205_ = 1'b1;
default : new_n3205_ = 1'b0;
endcase
casez ({new_n153_, new_n196_, new_n3418_})
3'b11? : new_n3206_ = 1'b1;
3'b??1 : new_n3206_ = 1'b1;
default : new_n3206_ = 1'b0;
endcase
casez ({new_n204_, new_n321_, new_n994_})
3'b11? : new_n3207_ = 1'b1;
3'b??1 : new_n3207_ = 1'b1;
default : new_n3207_ = 1'b0;
endcase
casez ({new_n313_, new_n2960_})
2'b00 : new_n3208_ = 1'b1;
default : new_n3208_ = 1'b0;
endcase
casez ({new_n139_, new_n208_, new_n3394_})
3'b11? : new_n3209_ = 1'b1;
3'b??1 : new_n3209_ = 1'b1;
default : new_n3209_ = 1'b0;
endcase
casez ({new_n177_, new_n2961_})
2'b00 : new_n3210_ = 1'b1;
default : new_n3210_ = 1'b0;
endcase
casez ({new_n153_, new_n2962_, new_n214_, new_n231_})
4'b11?? : new_n3211_ = 1'b1;
4'b??11 : new_n3211_ = 1'b1;
default : new_n3211_ = 1'b0;
endcase
casez ({y[2], new_n2963_, v[2], new_n180_})
4'b11?? : new_n3212_ = 1'b1;
4'b??11 : new_n3212_ = 1'b1;
default : new_n3212_ = 1'b0;
endcase
casez ({new_n342_, new_n2964_})
2'b00 : new_n3213_ = 1'b1;
default : new_n3213_ = 1'b0;
endcase
casez ({new_n3382_, new_n2966_})
2'b1? : new_n3214_ = 1'b1;
2'b?1 : new_n3214_ = 1'b1;
default : new_n3214_ = 1'b0;
endcase
casez ({new_n80_, new_n97_, new_n209_})
3'b01? : new_n3215_ = 1'b1;
3'b??1 : new_n3215_ = 1'b1;
default : new_n3215_ = 1'b0;
endcase
casez ({new_n187_, new_n210_})
2'b00 : new_n3216_ = 1'b1;
default : new_n3216_ = 1'b0;
endcase
casez ({y[0], new_n212_, new_n98_, new_n137_})
4'b11?? : new_n3217_ = 1'b1;
4'b??11 : new_n3217_ = 1'b1;
default : new_n3217_ = 1'b0;
endcase
casez ({new_n80_, new_n144_, new_n90_, new_n212_})
4'b11?? : new_n3218_ = 1'b1;
4'b??11 : new_n3218_ = 1'b1;
default : new_n3218_ = 1'b0;
endcase
casez ({new_n140_, new_n213_})
2'b00 : new_n3219_ = 1'b1;
default : new_n3219_ = 1'b0;
endcase
casez ({x[1], new_n184_, new_n87_, new_n385_})
4'b01?? : new_n3220_ = 1'b1;
4'b??11 : new_n3220_ = 1'b1;
default : new_n3220_ = 1'b0;
endcase
casez ({new_n79_, new_n83_, new_n214_})
3'b10? : new_n3221_ = 1'b1;
3'b??1 : new_n3221_ = 1'b1;
default : new_n3221_ = 1'b0;
endcase
casez ({new_n184_, new_n385_})
2'b00 : new_n3222_ = 1'b1;
default : new_n3222_ = 1'b0;
endcase
casez ({y[2], new_n79_, new_n214_})
3'b00? : new_n3223_ = 1'b1;
3'b??1 : new_n3223_ = 1'b1;
default : new_n3223_ = 1'b0;
endcase
casez ({new_n255_, new_n386_})
2'b00 : new_n3224_ = 1'b1;
default : new_n3224_ = 1'b0;
endcase
casez ({new_n207_, new_n386_, new_n216_, new_n306_})
4'b11?? : new_n3225_ = 1'b1;
4'b??11 : new_n3225_ = 1'b1;
default : new_n3225_ = 1'b0;
endcase
casez ({new_n170_, new_n215_})
2'b00 : new_n3226_ = 1'b1;
default : new_n3226_ = 1'b0;
endcase
casez ({new_n196_, new_n215_})
2'b00 : new_n3227_ = 1'b1;
default : new_n3227_ = 1'b0;
endcase
casez ({new_n123_, new_n215_, new_n3405_})
3'b11? : new_n3228_ = 1'b1;
3'b??1 : new_n3228_ = 1'b1;
default : new_n3228_ = 1'b0;
endcase
casez ({new_n151_, new_n215_})
2'b00 : new_n3229_ = 1'b1;
default : new_n3229_ = 1'b0;
endcase
casez ({new_n127_, new_n216_, new_n169_, new_n205_})
4'b11?? : new_n3230_ = 1'b1;
4'b??11 : new_n3230_ = 1'b1;
default : new_n3230_ = 1'b0;
endcase
casez ({new_n3529_, new_n145_})
2'b1? : new_n3231_ = 1'b1;
2'b?1 : new_n3231_ = 1'b1;
default : new_n3231_ = 1'b0;
endcase
casez ({new_n142_, new_n144_, new_n148_, new_n217_})
4'b11?? : new_n3232_ = 1'b1;
4'b??11 : new_n3232_ = 1'b1;
default : new_n3232_ = 1'b0;
endcase
casez ({new_n3504_, new_n3532_})
2'b1? : new_n3233_ = 1'b1;
2'b?1 : new_n3233_ = 1'b1;
default : new_n3233_ = 1'b0;
endcase
casez ({new_n198_, new_n219_})
2'b00 : new_n3234_ = 1'b1;
default : new_n3234_ = 1'b0;
endcase
casez ({new_n82_, new_n220_})
2'b00 : new_n3235_ = 1'b1;
default : new_n3235_ = 1'b0;
endcase
casez ({new_n190_, new_n210_, new_n191_, new_n220_})
4'b11?? : new_n3236_ = 1'b1;
4'b??11 : new_n3236_ = 1'b1;
default : new_n3236_ = 1'b0;
endcase
casez ({new_n3537_, new_n90_, new_n97_})
3'b1?? : new_n3237_ = 1'b1;
3'b?11 : new_n3237_ = 1'b1;
default : new_n3237_ = 1'b0;
endcase
casez ({new_n84_, new_n221_, new_n120_})
3'b01? : new_n3238_ = 1'b1;
3'b??1 : new_n3238_ = 1'b1;
default : new_n3238_ = 1'b0;
endcase
casez ({new_n95_, new_n221_})
2'b00 : new_n3239_ = 1'b1;
default : new_n3239_ = 1'b0;
endcase
casez ({new_n191_, new_n260_, new_n344_, new_n411_})
4'b11?? : new_n3240_ = 1'b1;
4'b??11 : new_n3240_ = 1'b1;
default : new_n3240_ = 1'b0;
endcase
casez ({new_n220_, new_n222_})
2'b00 : new_n3241_ = 1'b1;
default : new_n3241_ = 1'b0;
endcase
casez ({new_n161_, new_n411_, new_n230_, new_n241_})
4'b11?? : new_n3242_ = 1'b1;
4'b??11 : new_n3242_ = 1'b1;
default : new_n3242_ = 1'b0;
endcase
casez ({new_n187_, new_n706_, new_n210_, new_n231_})
4'b11?? : new_n3243_ = 1'b1;
4'b??11 : new_n3243_ = 1'b1;
default : new_n3243_ = 1'b0;
endcase
casez ({new_n189_, new_n411_, new_n209_, new_n239_})
4'b11?? : new_n3244_ = 1'b1;
4'b??11 : new_n3244_ = 1'b1;
default : new_n3244_ = 1'b0;
endcase
casez ({v[1], new_n222_, new_n3553_})
3'b11? : new_n3245_ = 1'b1;
3'b??1 : new_n3245_ = 1'b1;
default : new_n3245_ = 1'b0;
endcase
casez ({new_n158_, new_n213_, new_n177_, new_n222_})
4'b11?? : new_n3246_ = 1'b1;
4'b??11 : new_n3246_ = 1'b1;
default : new_n3246_ = 1'b0;
endcase
casez ({new_n170_, new_n222_, new_n201_, new_n213_})
4'b11?? : new_n3247_ = 1'b1;
4'b??11 : new_n3247_ = 1'b1;
default : new_n3247_ = 1'b0;
endcase
casez ({new_n94_, new_n99_, new_n222_})
3'b10? : new_n3248_ = 1'b1;
3'b??1 : new_n3248_ = 1'b1;
default : new_n3248_ = 1'b0;
endcase
casez ({new_n151_, new_n155_, new_n218_, new_n223_})
4'b11?? : new_n3249_ = 1'b1;
4'b??11 : new_n3249_ = 1'b1;
default : new_n3249_ = 1'b0;
endcase
casez ({new_n3545_, new_n3585_})
2'b1? : new_n3250_ = 1'b1;
2'b?1 : new_n3250_ = 1'b1;
default : new_n3250_ = 1'b0;
endcase
casez ({new_n96_, new_n190_, new_n155_, new_n224_})
4'b11?? : new_n3251_ = 1'b1;
4'b??11 : new_n3251_ = 1'b1;
default : new_n3251_ = 1'b0;
endcase
casez ({new_n159_, new_n417_, new_n3406_})
3'b11? : new_n3252_ = 1'b1;
3'b??1 : new_n3252_ = 1'b1;
default : new_n3252_ = 1'b0;
endcase
casez ({new_n79_, new_n224_, new_n3584_})
3'b11? : new_n3253_ = 1'b1;
3'b??1 : new_n3253_ = 1'b1;
default : new_n3253_ = 1'b0;
endcase
casez ({new_n144_, new_n226_})
2'b00 : new_n3254_ = 1'b1;
default : new_n3254_ = 1'b0;
endcase
casez ({new_n141_, new_n228_})
2'b00 : new_n3255_ = 1'b1;
default : new_n3255_ = 1'b0;
endcase
casez ({new_n115_, new_n127_, new_n214_, new_n228_})
4'b11?? : new_n3256_ = 1'b1;
4'b??11 : new_n3256_ = 1'b1;
default : new_n3256_ = 1'b0;
endcase
casez ({new_n118_, new_n120_})
2'b00 : new_n3257_ = 1'b1;
default : new_n3257_ = 1'b0;
endcase
casez ({new_n173_, new_n228_})
2'b00 : new_n3258_ = 1'b1;
default : new_n3258_ = 1'b0;
endcase
casez ({new_n83_, new_n427_, new_n84_, new_n285_})
4'b11?? : new_n3259_ = 1'b1;
4'b??11 : new_n3259_ = 1'b1;
default : new_n3259_ = 1'b0;
endcase
casez ({new_n183_, new_n229_})
2'b00 : new_n3260_ = 1'b1;
default : new_n3260_ = 1'b0;
endcase
casez ({new_n3497_, new_n167_, new_n427_})
3'b1?? : new_n3261_ = 1'b1;
3'b?11 : new_n3261_ = 1'b1;
default : new_n3261_ = 1'b0;
endcase
casez ({new_n196_, new_n229_})
2'b00 : new_n3262_ = 1'b1;
default : new_n3262_ = 1'b0;
endcase
casez ({new_n138_, new_n229_})
2'b00 : new_n3263_ = 1'b1;
default : new_n3263_ = 1'b0;
endcase
casez ({new_n194_, new_n432_})
2'b00 : new_n3264_ = 1'b1;
default : new_n3264_ = 1'b0;
endcase
casez ({new_n89_, new_n139_, new_n3437_})
3'b11? : new_n3265_ = 1'b1;
3'b??1 : new_n3265_ = 1'b1;
default : new_n3265_ = 1'b0;
endcase
casez ({x[2], new_n198_, u[1], new_n432_})
4'b11?? : new_n3266_ = 1'b1;
4'b??11 : new_n3266_ = 1'b1;
default : new_n3266_ = 1'b0;
endcase
casez ({new_n3422_, new_n3438_})
2'b1? : new_n3267_ = 1'b1;
2'b?1 : new_n3267_ = 1'b1;
default : new_n3267_ = 1'b0;
endcase
casez ({new_n3386_, new_n3438_})
2'b1? : new_n3268_ = 1'b1;
2'b?1 : new_n3268_ = 1'b1;
default : new_n3268_ = 1'b0;
endcase
casez ({new_n162_, new_n230_, new_n207_, new_n224_})
4'b11?? : new_n3269_ = 1'b1;
4'b??11 : new_n3269_ = 1'b1;
default : new_n3269_ = 1'b0;
endcase
casez ({new_n153_, new_n230_, new_n216_, new_n224_})
4'b11?? : new_n3270_ = 1'b1;
4'b??11 : new_n3270_ = 1'b1;
default : new_n3270_ = 1'b0;
endcase
casez ({new_n137_, new_n433_})
2'b00 : new_n3271_ = 1'b1;
default : new_n3271_ = 1'b0;
endcase
casez ({new_n151_, new_n230_})
2'b00 : new_n3272_ = 1'b1;
default : new_n3272_ = 1'b0;
endcase
casez ({x[2], new_n137_, new_n187_, new_n437_})
4'b01?? : new_n3273_ = 1'b1;
4'b??11 : new_n3273_ = 1'b1;
default : new_n3273_ = 1'b0;
endcase
casez ({new_n170_, new_n438_, new_n217_, new_n223_})
4'b11?? : new_n3274_ = 1'b1;
4'b??11 : new_n3274_ = 1'b1;
default : new_n3274_ = 1'b0;
endcase
casez ({new_n205_, new_n438_})
2'b00 : new_n3275_ = 1'b1;
default : new_n3275_ = 1'b0;
endcase
casez ({new_n123_, new_n231_})
2'b00 : new_n3276_ = 1'b1;
default : new_n3276_ = 1'b0;
endcase
casez ({new_n3506_, new_n94_, new_n728_})
3'b1?? : new_n3277_ = 1'b1;
3'b?11 : new_n3277_ = 1'b1;
default : new_n3277_ = 1'b0;
endcase
casez ({new_n190_, new_n728_, new_n217_, new_n264_})
4'b11?? : new_n3278_ = 1'b1;
4'b??11 : new_n3278_ = 1'b1;
default : new_n3278_ = 1'b0;
endcase
casez ({new_n138_, new_n260_, new_n469_, new_n730_})
4'b11?? : new_n3279_ = 1'b1;
4'b??11 : new_n3279_ = 1'b1;
default : new_n3279_ = 1'b0;
endcase
casez ({new_n177_, new_n234_})
2'b00 : new_n3280_ = 1'b1;
default : new_n3280_ = 1'b0;
endcase
casez ({new_n91_, new_n445_})
2'b00 : new_n3281_ = 1'b1;
default : new_n3281_ = 1'b0;
endcase
casez ({u[1], new_n92_, new_n1092_})
3'b01? : new_n3282_ = 1'b1;
3'b??1 : new_n3282_ = 1'b1;
default : new_n3282_ = 1'b0;
endcase
casez ({y[2], new_n152_, v[1], new_n1094_})
4'b11?? : new_n3283_ = 1'b1;
4'b??01 : new_n3283_ = 1'b1;
default : new_n3283_ = 1'b0;
endcase
casez ({new_n293_, new_n1095_})
2'b00 : new_n3284_ = 1'b1;
default : new_n3284_ = 1'b0;
endcase
casez ({new_n137_, new_n356_, new_n343_, new_n1096_})
4'b11?? : new_n3285_ = 1'b1;
4'b??11 : new_n3285_ = 1'b1;
default : new_n3285_ = 1'b0;
endcase
casez ({x[1], new_n1097_, new_n729_})
3'b01? : new_n3286_ = 1'b1;
3'b??1 : new_n3286_ = 1'b1;
default : new_n3286_ = 1'b0;
endcase
casez ({new_n153_, new_n1097_, new_n210_, new_n216_})
4'b11?? : new_n3287_ = 1'b1;
4'b??11 : new_n3287_ = 1'b1;
default : new_n3287_ = 1'b0;
endcase
casez ({new_n192_, new_n237_})
2'b00 : new_n3288_ = 1'b1;
default : new_n3288_ = 1'b0;
endcase
casez ({new_n190_, new_n1796_, new_n226_, new_n444_})
4'b11?? : new_n3289_ = 1'b1;
4'b??11 : new_n3289_ = 1'b1;
default : new_n3289_ = 1'b0;
endcase
casez ({new_n135_, new_n1797_})
2'b00 : new_n3290_ = 1'b1;
default : new_n3290_ = 1'b0;
endcase
casez ({new_n244_, new_n1798_})
2'b00 : new_n3291_ = 1'b1;
default : new_n3291_ = 1'b0;
endcase
casez ({new_n95_, new_n154_, new_n207_, new_n239_})
4'b11?? : new_n3292_ = 1'b1;
4'b??11 : new_n3292_ = 1'b1;
default : new_n3292_ = 1'b0;
endcase
casez ({new_n598_, new_n1802_})
2'b00 : new_n3293_ = 1'b1;
default : new_n3293_ = 1'b0;
endcase
casez ({u[0], new_n205_, new_n1805_})
3'b01? : new_n3294_ = 1'b1;
3'b??1 : new_n3294_ = 1'b1;
default : new_n3294_ = 1'b0;
endcase
casez ({new_n161_, new_n309_, new_n1806_})
3'b11? : new_n3295_ = 1'b1;
3'b??1 : new_n3295_ = 1'b1;
default : new_n3295_ = 1'b0;
endcase
casez ({new_n169_, new_n200_, new_n1806_})
3'b11? : new_n3296_ = 1'b1;
3'b??1 : new_n3296_ = 1'b1;
default : new_n3296_ = 1'b0;
endcase
casez ({new_n220_, new_n239_})
2'b00 : new_n3297_ = 1'b1;
default : new_n3297_ = 1'b0;
endcase
casez ({new_n89_, new_n127_, new_n1807_})
3'b01? : new_n3298_ = 1'b1;
3'b??1 : new_n3298_ = 1'b1;
default : new_n3298_ = 1'b0;
endcase
casez ({new_n198_, new_n241_})
2'b00 : new_n3299_ = 1'b1;
default : new_n3299_ = 1'b0;
endcase
casez ({new_n151_, new_n241_, new_n153_, new_n178_})
4'b11?? : new_n3300_ = 1'b1;
4'b??11 : new_n3300_ = 1'b1;
default : new_n3300_ = 1'b0;
endcase
casez ({new_n118_, new_n241_})
2'b00 : new_n3301_ = 1'b1;
default : new_n3301_ = 1'b0;
endcase
casez ({new_n167_, new_n198_, new_n211_, new_n242_})
4'b11?? : new_n3302_ = 1'b1;
4'b??11 : new_n3302_ = 1'b1;
default : new_n3302_ = 1'b0;
endcase
casez ({new_n201_, new_n242_})
2'b00 : new_n3303_ = 1'b1;
default : new_n3303_ = 1'b0;
endcase
casez ({new_n118_, new_n189_, new_n148_, new_n244_})
4'b11?? : new_n3304_ = 1'b1;
4'b??11 : new_n3304_ = 1'b1;
default : new_n3304_ = 1'b0;
endcase
casez ({new_n3540_, new_n215_, new_n244_})
3'b1?? : new_n3305_ = 1'b1;
3'b?11 : new_n3305_ = 1'b1;
default : new_n3305_ = 1'b0;
endcase
casez ({new_n129_, new_n273_, new_n145_, new_n469_})
4'b11?? : new_n3306_ = 1'b1;
4'b??11 : new_n3306_ = 1'b1;
default : new_n3306_ = 1'b0;
endcase
casez ({new_n215_, new_n247_, new_n220_, new_n229_})
4'b11?? : new_n3307_ = 1'b1;
4'b??11 : new_n3307_ = 1'b1;
default : new_n3307_ = 1'b0;
endcase
casez ({new_n223_, new_n248_})
2'b00 : new_n3308_ = 1'b1;
default : new_n3308_ = 1'b0;
endcase
casez ({new_n89_, new_n206_, new_n3562_})
3'b01? : new_n3309_ = 1'b1;
3'b??1 : new_n3309_ = 1'b1;
default : new_n3309_ = 1'b0;
endcase
casez ({new_n104_, new_n219_, new_n212_, new_n248_})
4'b11?? : new_n3310_ = 1'b1;
4'b??11 : new_n3310_ = 1'b1;
default : new_n3310_ = 1'b0;
endcase
casez ({new_n148_, new_n248_, new_n3424_})
3'b11? : new_n3311_ = 1'b1;
3'b??1 : new_n3311_ = 1'b1;
default : new_n3311_ = 1'b0;
endcase
casez ({new_n151_, new_n444_, new_n194_, new_n476_})
4'b11?? : new_n3312_ = 1'b1;
4'b??11 : new_n3312_ = 1'b1;
default : new_n3312_ = 1'b0;
endcase
casez ({v[0], new_n250_, new_n3453_})
3'b01? : new_n3313_ = 1'b1;
3'b??1 : new_n3313_ = 1'b1;
default : new_n3313_ = 1'b0;
endcase
casez ({new_n207_, new_n250_})
2'b00 : new_n3314_ = 1'b1;
default : new_n3314_ = 1'b0;
endcase
casez ({new_n118_, new_n250_})
2'b00 : new_n3315_ = 1'b1;
default : new_n3315_ = 1'b0;
endcase
casez ({new_n216_, new_n250_})
2'b00 : new_n3316_ = 1'b1;
default : new_n3316_ = 1'b0;
endcase
casez ({v[0], new_n77_})
2'b10 : new_n3317_ = 1'b1;
default : new_n3317_ = 1'b0;
endcase
casez ({new_n142_, new_n251_})
2'b11 : new_n3318_ = 1'b1;
default : new_n3318_ = 1'b0;
endcase
casez ({new_n115_, new_n765_})
2'b11 : new_n3319_ = 1'b1;
default : new_n3319_ = 1'b0;
endcase
casez ({new_n95_, new_n141_})
2'b01 : new_n3320_ = 1'b1;
default : new_n3320_ = 1'b0;
endcase
casez ({new_n139_, new_n254_})
2'b11 : new_n3321_ = 1'b1;
default : new_n3321_ = 1'b0;
endcase
casez ({x[1], new_n251_})
2'b01 : new_n3322_ = 1'b1;
default : new_n3322_ = 1'b0;
endcase
casez ({new_n169_, new_n255_})
2'b11 : new_n3323_ = 1'b1;
default : new_n3323_ = 1'b0;
endcase
casez ({new_n177_, new_n489_})
2'b11 : new_n3324_ = 1'b1;
default : new_n3324_ = 1'b0;
endcase
casez ({new_n242_, new_n489_})
2'b11 : new_n3325_ = 1'b1;
default : new_n3325_ = 1'b0;
endcase
casez ({new_n88_, new_n143_})
2'b01 : new_n3326_ = 1'b1;
default : new_n3326_ = 1'b0;
endcase
casez ({new_n191_, new_n257_})
2'b11 : new_n3327_ = 1'b1;
default : new_n3327_ = 1'b0;
endcase
casez ({new_n159_, new_n257_})
2'b11 : new_n3328_ = 1'b1;
default : new_n3328_ = 1'b0;
endcase
casez ({new_n207_, new_n258_})
2'b11 : new_n3329_ = 1'b1;
default : new_n3329_ = 1'b0;
endcase
casez ({new_n131_, new_n258_})
2'b11 : new_n3330_ = 1'b1;
default : new_n3330_ = 1'b0;
endcase
casez ({new_n182_, new_n260_})
2'b11 : new_n3331_ = 1'b1;
default : new_n3331_ = 1'b0;
endcase
casez ({new_n183_, new_n260_})
2'b11 : new_n3332_ = 1'b1;
default : new_n3332_ = 1'b0;
endcase
casez ({new_n200_, new_n260_})
2'b11 : new_n3333_ = 1'b1;
default : new_n3333_ = 1'b0;
endcase
casez ({new_n207_, new_n261_})
2'b11 : new_n3334_ = 1'b1;
default : new_n3334_ = 1'b0;
endcase
casez ({new_n85_, new_n508_})
2'b11 : new_n3335_ = 1'b1;
default : new_n3335_ = 1'b0;
endcase
casez ({new_n160_, new_n508_})
2'b11 : new_n3336_ = 1'b1;
default : new_n3336_ = 1'b0;
endcase
casez ({new_n160_, new_n264_})
2'b11 : new_n3337_ = 1'b1;
default : new_n3337_ = 1'b0;
endcase
casez ({new_n178_, new_n264_})
2'b11 : new_n3338_ = 1'b1;
default : new_n3338_ = 1'b0;
endcase
casez ({new_n159_, new_n509_})
2'b11 : new_n3339_ = 1'b1;
default : new_n3339_ = 1'b0;
endcase
casez ({new_n237_, new_n264_})
2'b11 : new_n3340_ = 1'b1;
default : new_n3340_ = 1'b0;
endcase
casez ({new_n139_, new_n266_})
2'b11 : new_n3341_ = 1'b1;
default : new_n3341_ = 1'b0;
endcase
casez ({new_n101_, new_n152_})
2'b11 : new_n3342_ = 1'b1;
default : new_n3342_ = 1'b0;
endcase
casez ({new_n177_, new_n531_})
2'b11 : new_n3343_ = 1'b1;
default : new_n3343_ = 1'b0;
endcase
casez ({new_n160_, new_n531_})
2'b11 : new_n3344_ = 1'b1;
default : new_n3344_ = 1'b0;
endcase
casez ({new_n194_, new_n532_})
2'b11 : new_n3345_ = 1'b1;
default : new_n3345_ = 1'b0;
endcase
casez ({new_n97_, new_n532_})
2'b11 : new_n3346_ = 1'b1;
default : new_n3346_ = 1'b0;
endcase
casez ({new_n87_, new_n156_})
2'b11 : new_n3347_ = 1'b1;
default : new_n3347_ = 1'b0;
endcase
casez ({new_n82_, new_n274_})
2'b01 : new_n3348_ = 1'b1;
default : new_n3348_ = 1'b0;
endcase
casez ({new_n145_, new_n274_})
2'b11 : new_n3349_ = 1'b1;
default : new_n3349_ = 1'b0;
endcase
casez ({new_n177_, new_n274_})
2'b11 : new_n3350_ = 1'b1;
default : new_n3350_ = 1'b0;
endcase
casez ({new_n148_, new_n158_})
2'b11 : new_n3351_ = 1'b1;
default : new_n3351_ = 1'b0;
endcase
casez ({new_n161_, new_n274_})
2'b11 : new_n3352_ = 1'b1;
default : new_n3352_ = 1'b0;
endcase
casez ({new_n97_, new_n822_})
2'b11 : new_n3353_ = 1'b1;
default : new_n3353_ = 1'b0;
endcase
casez ({new_n261_, new_n284_})
2'b11 : new_n3354_ = 1'b1;
default : new_n3354_ = 1'b0;
endcase
casez ({new_n123_, new_n162_})
2'b11 : new_n3355_ = 1'b1;
default : new_n3355_ = 1'b0;
endcase
casez ({new_n150_, new_n285_})
2'b11 : new_n3356_ = 1'b1;
default : new_n3356_ = 1'b0;
endcase
casez ({new_n94_, new_n165_})
2'b01 : new_n3357_ = 1'b1;
default : new_n3357_ = 1'b0;
endcase
casez ({new_n231_, new_n287_})
2'b11 : new_n3358_ = 1'b1;
default : new_n3358_ = 1'b0;
endcase
casez ({new_n205_, new_n287_})
2'b11 : new_n3359_ = 1'b1;
default : new_n3359_ = 1'b0;
endcase
casez ({new_n87_, new_n565_})
2'b01 : new_n3360_ = 1'b1;
default : new_n3360_ = 1'b0;
endcase
casez ({new_n80_, new_n167_})
2'b01 : new_n3361_ = 1'b1;
default : new_n3361_ = 1'b0;
endcase
casez ({new_n95_, new_n169_})
2'b11 : new_n3362_ = 1'b1;
default : new_n3362_ = 1'b0;
endcase
casez ({u[2], new_n293_})
2'b01 : new_n3363_ = 1'b1;
default : new_n3363_ = 1'b0;
endcase
casez ({x[1], new_n170_})
2'b01 : new_n3364_ = 1'b1;
default : new_n3364_ = 1'b0;
endcase
casez ({new_n129_, new_n305_})
2'b11 : new_n3365_ = 1'b1;
default : new_n3365_ = 1'b0;
endcase
casez ({new_n150_, new_n305_})
2'b11 : new_n3366_ = 1'b1;
default : new_n3366_ = 1'b0;
endcase
casez ({new_n131_, new_n174_})
2'b11 : new_n3367_ = 1'b1;
default : new_n3367_ = 1'b0;
endcase
casez ({new_n153_, new_n301_})
2'b11 : new_n3368_ = 1'b1;
default : new_n3368_ = 1'b0;
endcase
casez ({new_n274_, new_n301_})
2'b11 : new_n3369_ = 1'b1;
default : new_n3369_ = 1'b0;
endcase
casez ({new_n198_, new_n307_})
2'b11 : new_n3370_ = 1'b1;
default : new_n3370_ = 1'b0;
endcase
casez ({new_n126_, new_n599_})
2'b11 : new_n3371_ = 1'b1;
default : new_n3371_ = 1'b0;
endcase
casez ({new_n199_, new_n313_})
2'b11 : new_n3372_ = 1'b1;
default : new_n3372_ = 1'b0;
endcase
casez ({new_n182_, new_n316_})
2'b11 : new_n3373_ = 1'b1;
default : new_n3373_ = 1'b0;
endcase
casez ({new_n183_, new_n316_})
2'b11 : new_n3374_ = 1'b1;
default : new_n3374_ = 1'b0;
endcase
casez ({x[2], new_n316_})
2'b11 : new_n3375_ = 1'b1;
default : new_n3375_ = 1'b0;
endcase
casez ({new_n103_, new_n317_})
2'b11 : new_n3376_ = 1'b1;
default : new_n3376_ = 1'b0;
endcase
casez ({new_n151_, new_n316_})
2'b11 : new_n3377_ = 1'b1;
default : new_n3377_ = 1'b0;
endcase
casez ({new_n96_, new_n2509_})
2'b11 : new_n3378_ = 1'b1;
default : new_n3378_ = 1'b0;
endcase
casez ({new_n184_, new_n321_})
2'b11 : new_n3379_ = 1'b1;
default : new_n3379_ = 1'b0;
endcase
casez ({new_n95_, new_n321_})
2'b11 : new_n3380_ = 1'b1;
default : new_n3380_ = 1'b0;
endcase
casez ({new_n96_, new_n615_})
2'b10 : new_n3381_ = 1'b1;
default : new_n3381_ = 1'b0;
endcase
casez ({x[2], new_n616_})
2'b11 : new_n3382_ = 1'b1;
default : new_n3382_ = 1'b0;
endcase
casez ({new_n189_, new_n332_})
2'b11 : new_n3383_ = 1'b1;
default : new_n3383_ = 1'b0;
endcase
casez ({v[1], new_n190_})
2'b11 : new_n3384_ = 1'b1;
default : new_n3384_ = 1'b0;
endcase
casez ({new_n305_, new_n338_})
2'b11 : new_n3385_ = 1'b1;
default : new_n3385_ = 1'b0;
endcase
casez ({new_n187_, new_n338_})
2'b11 : new_n3386_ = 1'b1;
default : new_n3386_ = 1'b0;
endcase
casez ({new_n145_, new_n194_})
2'b11 : new_n3387_ = 1'b1;
default : new_n3387_ = 1'b0;
endcase
casez ({new_n184_, new_n194_})
2'b11 : new_n3388_ = 1'b1;
default : new_n3388_ = 1'b0;
endcase
casez ({new_n77_, new_n99_})
2'b01 : new_n3389_ = 1'b1;
default : new_n3389_ = 1'b0;
endcase
casez ({new_n170_, new_n343_})
2'b11 : new_n3390_ = 1'b1;
default : new_n3390_ = 1'b0;
endcase
casez ({new_n321_, new_n344_})
2'b11 : new_n3391_ = 1'b1;
default : new_n3391_ = 1'b0;
endcase
casez ({new_n127_, new_n344_})
2'b11 : new_n3392_ = 1'b1;
default : new_n3392_ = 1'b0;
endcase
casez ({new_n220_, new_n346_})
2'b11 : new_n3393_ = 1'b1;
default : new_n3393_ = 1'b0;
endcase
casez ({new_n183_, new_n198_})
2'b11 : new_n3394_ = 1'b1;
default : new_n3394_ = 1'b0;
endcase
casez ({new_n178_, new_n198_})
2'b11 : new_n3395_ = 1'b1;
default : new_n3395_ = 1'b0;
endcase
casez ({new_n127_, new_n347_})
2'b11 : new_n3396_ = 1'b1;
default : new_n3396_ = 1'b0;
endcase
casez ({new_n94_, new_n347_})
2'b11 : new_n3397_ = 1'b1;
default : new_n3397_ = 1'b0;
endcase
casez ({new_n77_, new_n100_})
2'b11 : new_n3398_ = 1'b1;
default : new_n3398_ = 1'b0;
endcase
casez ({new_n115_, new_n201_})
2'b11 : new_n3399_ = 1'b1;
default : new_n3399_ = 1'b0;
endcase
casez ({new_n118_, new_n201_})
2'b11 : new_n3400_ = 1'b1;
default : new_n3400_ = 1'b0;
endcase
casez ({new_n151_, new_n358_})
2'b11 : new_n3401_ = 1'b1;
default : new_n3401_ = 1'b0;
endcase
casez ({new_n182_, new_n356_})
2'b11 : new_n3402_ = 1'b1;
default : new_n3402_ = 1'b0;
endcase
casez ({new_n118_, new_n204_})
2'b11 : new_n3403_ = 1'b1;
default : new_n3403_ = 1'b0;
endcase
casez ({new_n189_, new_n204_})
2'b11 : new_n3404_ = 1'b1;
default : new_n3404_ = 1'b0;
endcase
casez ({new_n173_, new_n204_})
2'b11 : new_n3405_ = 1'b1;
default : new_n3405_ = 1'b0;
endcase
casez ({new_n160_, new_n358_})
2'b11 : new_n3406_ = 1'b1;
default : new_n3406_ = 1'b0;
endcase
casez ({new_n183_, new_n205_})
2'b11 : new_n3407_ = 1'b1;
default : new_n3407_ = 1'b0;
endcase
casez ({new_n145_, new_n363_})
2'b11 : new_n3408_ = 1'b1;
default : new_n3408_ = 1'b0;
endcase
casez ({new_n154_, new_n205_})
2'b11 : new_n3409_ = 1'b1;
default : new_n3409_ = 1'b0;
endcase
casez ({new_n200_, new_n205_})
2'b11 : new_n3410_ = 1'b1;
default : new_n3410_ = 1'b0;
endcase
casez ({new_n189_, new_n363_})
2'b11 : new_n3411_ = 1'b1;
default : new_n3411_ = 1'b0;
endcase
casez ({new_n147_, new_n654_})
2'b11 : new_n3412_ = 1'b1;
default : new_n3412_ = 1'b0;
endcase
casez ({new_n176_, new_n207_})
2'b11 : new_n3413_ = 1'b1;
default : new_n3413_ = 1'b0;
endcase
casez ({new_n182_, new_n207_})
2'b11 : new_n3414_ = 1'b1;
default : new_n3414_ = 1'b0;
endcase
casez ({new_n156_, new_n2914_})
2'b11 : new_n3415_ = 1'b1;
default : new_n3415_ = 1'b0;
endcase
casez ({v[0], new_n994_})
2'b01 : new_n3416_ = 1'b1;
default : new_n3416_ = 1'b0;
endcase
casez ({new_n200_, new_n369_})
2'b11 : new_n3417_ = 1'b1;
default : new_n3417_ = 1'b0;
endcase
casez ({new_n206_, new_n991_})
2'b11 : new_n3418_ = 1'b1;
default : new_n3418_ = 1'b0;
endcase
casez ({new_n357_, new_n2976_})
2'b11 : new_n3419_ = 1'b1;
default : new_n3419_ = 1'b0;
endcase
casez ({new_n151_, new_n211_})
2'b11 : new_n3420_ = 1'b1;
default : new_n3420_ = 1'b0;
endcase
casez ({new_n167_, new_n211_})
2'b11 : new_n3421_ = 1'b1;
default : new_n3421_ = 1'b0;
endcase
casez ({new_n184_, new_n211_})
2'b11 : new_n3422_ = 1'b1;
default : new_n3422_ = 1'b0;
endcase
casez ({new_n97_, new_n213_})
2'b01 : new_n3423_ = 1'b1;
default : new_n3423_ = 1'b0;
endcase
casez ({new_n182_, new_n212_})
2'b11 : new_n3424_ = 1'b1;
default : new_n3424_ = 1'b0;
endcase
casez ({new_n155_, new_n216_})
2'b11 : new_n3425_ = 1'b1;
default : new_n3425_ = 1'b0;
endcase
casez ({new_n184_, new_n216_})
2'b11 : new_n3426_ = 1'b1;
default : new_n3426_ = 1'b0;
endcase
casez ({new_n211_, new_n218_})
2'b11 : new_n3427_ = 1'b1;
default : new_n3427_ = 1'b0;
endcase
casez ({new_n184_, new_n219_})
2'b11 : new_n3428_ = 1'b1;
default : new_n3428_ = 1'b0;
endcase
casez ({new_n129_, new_n216_})
2'b11 : new_n3429_ = 1'b1;
default : new_n3429_ = 1'b0;
endcase
casez ({new_n192_, new_n222_})
2'b11 : new_n3430_ = 1'b1;
default : new_n3430_ = 1'b0;
endcase
casez ({new_n144_, new_n411_})
2'b11 : new_n3431_ = 1'b1;
default : new_n3431_ = 1'b0;
endcase
casez ({new_n153_, new_n222_})
2'b11 : new_n3432_ = 1'b1;
default : new_n3432_ = 1'b0;
endcase
casez ({new_n123_, new_n223_})
2'b11 : new_n3433_ = 1'b1;
default : new_n3433_ = 1'b0;
endcase
casez ({x[1], new_n223_})
2'b11 : new_n3434_ = 1'b1;
default : new_n3434_ = 1'b0;
endcase
casez ({new_n83_, new_n228_})
2'b01 : new_n3435_ = 1'b1;
default : new_n3435_ = 1'b0;
endcase
casez ({new_n199_, new_n432_})
2'b11 : new_n3436_ = 1'b1;
default : new_n3436_ = 1'b0;
endcase
casez ({new_n187_, new_n432_})
2'b11 : new_n3437_ = 1'b1;
default : new_n3437_ = 1'b0;
endcase
casez ({new_n301_, new_n432_})
2'b11 : new_n3438_ = 1'b1;
default : new_n3438_ = 1'b0;
endcase
casez ({new_n214_, new_n235_})
2'b11 : new_n3439_ = 1'b1;
default : new_n3439_ = 1'b0;
endcase
casez ({new_n84_, new_n235_})
2'b01 : new_n3440_ = 1'b1;
default : new_n3440_ = 1'b0;
endcase
casez ({new_n89_, new_n445_})
2'b11 : new_n3441_ = 1'b1;
default : new_n3441_ = 1'b0;
endcase
casez ({new_n423_, new_n3441_, new_n952_, new_n1343_})
4'b11?? : new_n3442_ = 1'b1;
4'b??11 : new_n3442_ = 1'b1;
default : new_n3442_ = 1'b0;
endcase
casez ({new_n97_, new_n1094_})
2'b11 : new_n3443_ = 1'b1;
default : new_n3443_ = 1'b0;
endcase
casez ({new_n154_, new_n1801_})
2'b11 : new_n3444_ = 1'b1;
default : new_n3444_ = 1'b0;
endcase
casez ({new_n100_, new_n1808_})
2'b01 : new_n3445_ = 1'b1;
default : new_n3445_ = 1'b0;
endcase
casez ({new_n174_, new_n241_})
2'b11 : new_n3446_ = 1'b1;
default : new_n3446_ = 1'b0;
endcase
casez ({new_n107_, new_n242_})
2'b01 : new_n3447_ = 1'b1;
default : new_n3447_ = 1'b0;
endcase
casez ({new_n209_, new_n242_})
2'b11 : new_n3448_ = 1'b1;
default : new_n3448_ = 1'b0;
endcase
casez ({new_n154_, new_n244_})
2'b11 : new_n3449_ = 1'b1;
default : new_n3449_ = 1'b0;
endcase
casez ({new_n88_, new_n135_})
2'b01 : new_n3450_ = 1'b1;
default : new_n3450_ = 1'b0;
endcase
casez ({x[2], new_n469_})
2'b01 : new_n3451_ = 1'b1;
default : new_n3451_ = 1'b0;
endcase
casez ({new_n131_, new_n248_})
2'b11 : new_n3452_ = 1'b1;
default : new_n3452_ = 1'b0;
endcase
casez ({new_n219_, new_n247_})
2'b11 : new_n3453_ = 1'b1;
default : new_n3453_ = 1'b0;
endcase
casez ({new_n247_, new_n249_})
2'b11 : new_n3454_ = 1'b1;
default : new_n3454_ = 1'b0;
endcase
casez ({new_n80_, new_n254_})
2'b01 : new_n3455_ = 1'b1;
default : new_n3455_ = 1'b0;
endcase
casez ({new_n89_, new_n143_})
2'b01 : new_n3456_ = 1'b1;
default : new_n3456_ = 1'b0;
endcase
casez ({new_n215_, new_n257_})
2'b11 : new_n3457_ = 1'b1;
default : new_n3457_ = 1'b0;
endcase
casez ({u[2], new_n258_})
2'b01 : new_n3458_ = 1'b1;
default : new_n3458_ = 1'b0;
endcase
casez ({new_n208_, new_n260_})
2'b11 : new_n3459_ = 1'b1;
default : new_n3459_ = 1'b0;
endcase
casez ({new_n201_, new_n260_})
2'b11 : new_n3460_ = 1'b1;
default : new_n3460_ = 1'b0;
endcase
casez ({u[1], new_n148_})
2'b11 : new_n3461_ = 1'b1;
default : new_n3461_ = 1'b0;
endcase
casez ({new_n204_, new_n264_})
2'b11 : new_n3462_ = 1'b1;
default : new_n3462_ = 1'b0;
endcase
casez ({new_n210_, new_n264_})
2'b11 : new_n3463_ = 1'b1;
default : new_n3463_ = 1'b0;
endcase
casez ({u[2], new_n151_})
2'b11 : new_n3464_ = 1'b1;
default : new_n3464_ = 1'b0;
endcase
casez ({u[1], new_n153_})
2'b01 : new_n3465_ = 1'b1;
default : new_n3465_ = 1'b0;
endcase
casez ({new_n153_, new_n155_})
2'b11 : new_n3466_ = 1'b1;
default : new_n3466_ = 1'b0;
endcase
casez ({v[1], new_n155_})
2'b01 : new_n3467_ = 1'b1;
default : new_n3467_ = 1'b0;
endcase
casez ({new_n167_, new_n275_})
2'b11 : new_n3468_ = 1'b1;
default : new_n3468_ = 1'b0;
endcase
casez ({new_n107_, new_n158_})
2'b01 : new_n3469_ = 1'b1;
default : new_n3469_ = 1'b0;
endcase
casez ({new_n127_, new_n158_})
2'b11 : new_n3470_ = 1'b1;
default : new_n3470_ = 1'b0;
endcase
casez ({y[2], new_n279_})
2'b01 : new_n3471_ = 1'b1;
default : new_n3471_ = 1'b0;
endcase
casez ({new_n92_, new_n160_})
2'b11 : new_n3472_ = 1'b1;
default : new_n3472_ = 1'b0;
endcase
casez ({new_n89_, new_n279_})
2'b11 : new_n3473_ = 1'b1;
default : new_n3473_ = 1'b0;
endcase
casez ({new_n115_, new_n159_})
2'b11 : new_n3474_ = 1'b1;
default : new_n3474_ = 1'b0;
endcase
casez ({new_n153_, new_n161_})
2'b11 : new_n3475_ = 1'b1;
default : new_n3475_ = 1'b0;
endcase
casez ({new_n153_, new_n285_})
2'b11 : new_n3476_ = 1'b1;
default : new_n3476_ = 1'b0;
endcase
casez ({x[1], new_n166_})
2'b01 : new_n3477_ = 1'b1;
default : new_n3477_ = 1'b0;
endcase
casez ({u[2], new_n167_})
2'b01 : new_n3478_ = 1'b1;
default : new_n3478_ = 1'b0;
endcase
casez ({new_n79_, new_n170_})
2'b11 : new_n3479_ = 1'b1;
default : new_n3479_ = 1'b0;
endcase
casez ({new_n83_, new_n299_})
2'b11 : new_n3480_ = 1'b1;
default : new_n3480_ = 1'b0;
endcase
casez ({new_n104_, new_n173_})
2'b11 : new_n3481_ = 1'b1;
default : new_n3481_ = 1'b0;
endcase
casez ({new_n84_, new_n173_})
2'b11 : new_n3482_ = 1'b1;
default : new_n3482_ = 1'b0;
endcase
casez ({new_n92_, new_n174_})
2'b11 : new_n3483_ = 1'b1;
default : new_n3483_ = 1'b0;
endcase
casez ({new_n118_, new_n174_})
2'b11 : new_n3484_ = 1'b1;
default : new_n3484_ = 1'b0;
endcase
casez ({new_n154_, new_n174_})
2'b11 : new_n3485_ = 1'b1;
default : new_n3485_ = 1'b0;
endcase
casez ({new_n115_, new_n307_})
2'b11 : new_n3486_ = 1'b1;
default : new_n3486_ = 1'b0;
endcase
casez ({new_n142_, new_n176_})
2'b11 : new_n3487_ = 1'b1;
default : new_n3487_ = 1'b0;
endcase
casez ({new_n162_, new_n176_})
2'b11 : new_n3488_ = 1'b1;
default : new_n3488_ = 1'b0;
endcase
casez ({new_n107_, new_n177_})
2'b01 : new_n3489_ = 1'b1;
default : new_n3489_ = 1'b0;
endcase
casez ({new_n139_, new_n173_})
2'b11 : new_n3490_ = 1'b1;
default : new_n3490_ = 1'b0;
endcase
casez ({new_n109_, new_n178_})
2'b01 : new_n3491_ = 1'b1;
default : new_n3491_ = 1'b0;
endcase
casez ({x[1], new_n178_})
2'b11 : new_n3492_ = 1'b1;
default : new_n3492_ = 1'b0;
endcase
casez ({y[2], new_n313_})
2'b11 : new_n3493_ = 1'b1;
default : new_n3493_ = 1'b0;
endcase
casez ({new_n148_, new_n315_})
2'b11 : new_n3494_ = 1'b1;
default : new_n3494_ = 1'b0;
endcase
casez ({new_n84_, new_n318_})
2'b11 : new_n3495_ = 1'b1;
default : new_n3495_ = 1'b0;
endcase
casez ({new_n89_, new_n318_})
2'b11 : new_n3496_ = 1'b1;
default : new_n3496_ = 1'b0;
endcase
casez ({new_n81_, new_n182_})
2'b11 : new_n3497_ = 1'b1;
default : new_n3497_ = 1'b0;
endcase
casez ({new_n82_, new_n182_})
2'b11 : new_n3498_ = 1'b1;
default : new_n3498_ = 1'b0;
endcase
casez ({new_n145_, new_n321_})
2'b11 : new_n3499_ = 1'b1;
default : new_n3499_ = 1'b0;
endcase
casez ({new_n142_, new_n187_})
2'b11 : new_n3500_ = 1'b1;
default : new_n3500_ = 1'b0;
endcase
casez ({new_n118_, new_n187_})
2'b11 : new_n3501_ = 1'b1;
default : new_n3501_ = 1'b0;
endcase
casez ({new_n153_, new_n189_})
2'b11 : new_n3502_ = 1'b1;
default : new_n3502_ = 1'b0;
endcase
casez ({y[2], new_n190_})
2'b11 : new_n3503_ = 1'b1;
default : new_n3503_ = 1'b0;
endcase
casez ({x[0], new_n190_})
2'b01 : new_n3504_ = 1'b1;
default : new_n3504_ = 1'b0;
endcase
casez ({new_n161_, new_n194_})
2'b11 : new_n3505_ = 1'b1;
default : new_n3505_ = 1'b0;
endcase
casez ({new_n84_, new_n342_})
2'b11 : new_n3506_ = 1'b1;
default : new_n3506_ = 1'b0;
endcase
casez ({x[1], new_n196_})
2'b11 : new_n3507_ = 1'b1;
default : new_n3507_ = 1'b0;
endcase
casez ({new_n95_, new_n343_})
2'b11 : new_n3508_ = 1'b1;
default : new_n3508_ = 1'b0;
endcase
casez ({new_n158_, new_n198_})
2'b11 : new_n3509_ = 1'b1;
default : new_n3509_ = 1'b0;
endcase
casez ({new_n77_, new_n198_})
2'b11 : new_n3510_ = 1'b1;
default : new_n3510_ = 1'b0;
endcase
casez ({u[2], new_n199_})
2'b11 : new_n3511_ = 1'b1;
default : new_n3511_ = 1'b0;
endcase
casez ({new_n109_, new_n200_})
2'b01 : new_n3512_ = 1'b1;
default : new_n3512_ = 1'b0;
endcase
casez ({new_n198_, new_n200_})
2'b11 : new_n3513_ = 1'b1;
default : new_n3513_ = 1'b0;
endcase
casez ({new_n115_, new_n200_})
2'b11 : new_n3514_ = 1'b1;
default : new_n3514_ = 1'b0;
endcase
casez ({x[1], new_n201_})
2'b01 : new_n3515_ = 1'b1;
default : new_n3515_ = 1'b0;
endcase
casez ({new_n159_, new_n209_})
2'b11 : new_n3516_ = 1'b1;
default : new_n3516_ = 1'b0;
endcase
casez ({new_n191_, new_n209_})
2'b11 : new_n3517_ = 1'b1;
default : new_n3517_ = 1'b0;
endcase
casez ({new_n187_, new_n209_})
2'b11 : new_n3518_ = 1'b1;
default : new_n3518_ = 1'b0;
endcase
casez ({new_n80_, new_n210_})
2'b11 : new_n3519_ = 1'b1;
default : new_n3519_ = 1'b0;
endcase
casez ({u[1], new_n211_})
2'b01 : new_n3520_ = 1'b1;
default : new_n3520_ = 1'b0;
endcase
casez ({u[1], new_n212_})
2'b11 : new_n3521_ = 1'b1;
default : new_n3521_ = 1'b0;
endcase
casez ({x[2], new_n212_})
2'b11 : new_n3522_ = 1'b1;
default : new_n3522_ = 1'b0;
endcase
casez ({new_n153_, new_n213_})
2'b11 : new_n3523_ = 1'b1;
default : new_n3523_ = 1'b0;
endcase
casez ({new_n140_, new_n214_})
2'b11 : new_n3524_ = 1'b1;
default : new_n3524_ = 1'b0;
endcase
casez ({new_n162_, new_n386_})
2'b11 : new_n3525_ = 1'b1;
default : new_n3525_ = 1'b0;
endcase
casez ({new_n123_, new_n363_})
2'b11 : new_n3526_ = 1'b1;
default : new_n3526_ = 1'b0;
endcase
casez ({new_n94_, new_n215_})
2'b11 : new_n3527_ = 1'b1;
default : new_n3527_ = 1'b0;
endcase
casez ({new_n159_, new_n216_})
2'b11 : new_n3528_ = 1'b1;
default : new_n3528_ = 1'b0;
endcase
casez ({y[2], new_n217_})
2'b01 : new_n3529_ = 1'b1;
default : new_n3529_ = 1'b0;
endcase
casez ({new_n100_, new_n216_})
2'b11 : new_n3530_ = 1'b1;
default : new_n3530_ = 1'b0;
endcase
casez ({new_n118_, new_n218_})
2'b11 : new_n3531_ = 1'b1;
default : new_n3531_ = 1'b0;
endcase
casez ({new_n88_, new_n218_})
2'b11 : new_n3532_ = 1'b1;
default : new_n3532_ = 1'b0;
endcase
casez ({new_n174_, new_n219_})
2'b11 : new_n3533_ = 1'b1;
default : new_n3533_ = 1'b0;
endcase
casez ({new_n86_, new_n219_})
2'b11 : new_n3534_ = 1'b1;
default : new_n3534_ = 1'b0;
endcase
casez ({u[1], new_n219_})
2'b11 : new_n3535_ = 1'b1;
default : new_n3535_ = 1'b0;
endcase
casez ({v[2], new_n219_})
2'b01 : new_n3536_ = 1'b1;
default : new_n3536_ = 1'b0;
endcase
casez ({v[1], new_n220_})
2'b01 : new_n3537_ = 1'b1;
default : new_n3537_ = 1'b0;
endcase
casez ({new_n97_, new_n221_})
2'b11 : new_n3538_ = 1'b1;
default : new_n3538_ = 1'b0;
endcase
casez ({x[0], new_n221_})
2'b01 : new_n3539_ = 1'b1;
default : new_n3539_ = 1'b0;
endcase
casez ({new_n160_, new_n221_})
2'b11 : new_n3540_ = 1'b1;
default : new_n3540_ = 1'b0;
endcase
casez ({u[1], new_n115_})
2'b11 : new_n3541_ = 1'b1;
default : new_n3541_ = 1'b0;
endcase
casez ({y[2], new_n222_})
2'b11 : new_n3542_ = 1'b1;
default : new_n3542_ = 1'b0;
endcase
casez ({new_n98_, new_n222_})
2'b11 : new_n3543_ = 1'b1;
default : new_n3543_ = 1'b0;
endcase
casez ({v[1], new_n116_})
2'b11 : new_n3544_ = 1'b1;
default : new_n3544_ = 1'b0;
endcase
casez ({u[2], new_n223_})
2'b01 : new_n3545_ = 1'b1;
default : new_n3545_ = 1'b0;
endcase
casez ({new_n139_, new_n224_})
2'b11 : new_n3546_ = 1'b1;
default : new_n3546_ = 1'b0;
endcase
casez ({new_n84_, new_n226_})
2'b11 : new_n3547_ = 1'b1;
default : new_n3547_ = 1'b0;
endcase
casez ({new_n97_, new_n228_})
2'b11 : new_n3548_ = 1'b1;
default : new_n3548_ = 1'b0;
endcase
casez ({new_n118_, new_n229_})
2'b11 : new_n3549_ = 1'b1;
default : new_n3549_ = 1'b0;
endcase
casez ({new_n131_, new_n230_})
2'b11 : new_n3550_ = 1'b1;
default : new_n3550_ = 1'b0;
endcase
casez ({new_n103_, new_n231_})
2'b11 : new_n3551_ = 1'b1;
default : new_n3551_ = 1'b0;
endcase
casez ({new_n98_, new_n235_})
2'b11 : new_n3552_ = 1'b1;
default : new_n3552_ = 1'b0;
endcase
casez ({new_n84_, new_n127_})
2'b01 : new_n3553_ = 1'b1;
default : new_n3553_ = 1'b0;
endcase
casez ({new_n95_, new_n238_})
2'b11 : new_n3554_ = 1'b1;
default : new_n3554_ = 1'b0;
endcase
casez ({new_n83_, new_n238_})
2'b11 : new_n3555_ = 1'b1;
default : new_n3555_ = 1'b0;
endcase
casez ({new_n178_, new_n241_})
2'b11 : new_n3556_ = 1'b1;
default : new_n3556_ = 1'b0;
endcase
casez ({new_n96_, new_n244_})
2'b11 : new_n3557_ = 1'b1;
default : new_n3557_ = 1'b0;
endcase
casez ({new_n79_, new_n133_})
2'b01 : new_n3558_ = 1'b1;
default : new_n3558_ = 1'b0;
endcase
casez ({new_n98_, new_n247_})
2'b11 : new_n3559_ = 1'b1;
default : new_n3559_ = 1'b0;
endcase
casez ({new_n109_, new_n248_})
2'b01 : new_n3560_ = 1'b1;
default : new_n3560_ = 1'b0;
endcase
casez ({new_n94_, new_n248_})
2'b11 : new_n3561_ = 1'b1;
default : new_n3561_ = 1'b0;
endcase
casez ({new_n198_, new_n248_})
2'b11 : new_n3562_ = 1'b1;
default : new_n3562_ = 1'b0;
endcase
casez ({new_n104_, new_n140_})
2'b11 : new_n3563_ = 1'b1;
default : new_n3563_ = 1'b0;
endcase
casez ({v[1], new_n143_})
2'b01 : new_n3564_ = 1'b1;
default : new_n3564_ = 1'b0;
endcase
casez ({y[2], new_n143_})
2'b01 : new_n3565_ = 1'b1;
default : new_n3565_ = 1'b0;
endcase
casez ({y[2], new_n143_})
2'b11 : new_n3566_ = 1'b1;
default : new_n3566_ = 1'b0;
endcase
casez ({new_n84_, new_n144_})
2'b11 : new_n3567_ = 1'b1;
default : new_n3567_ = 1'b0;
endcase
casez ({new_n88_, new_n145_})
2'b11 : new_n3568_ = 1'b1;
default : new_n3568_ = 1'b0;
endcase
casez ({new_n97_, new_n145_})
2'b11 : new_n3569_ = 1'b1;
default : new_n3569_ = 1'b0;
endcase
casez ({new_n85_, new_n148_})
2'b11 : new_n3570_ = 1'b1;
default : new_n3570_ = 1'b0;
endcase
casez ({x[2], new_n148_})
2'b01 : new_n3571_ = 1'b1;
default : new_n3571_ = 1'b0;
endcase
casez ({new_n90_, new_n148_})
2'b11 : new_n3572_ = 1'b1;
default : new_n3572_ = 1'b0;
endcase
casez ({new_n86_, new_n148_})
2'b11 : new_n3573_ = 1'b1;
default : new_n3573_ = 1'b0;
endcase
casez ({new_n92_, new_n151_})
2'b11 : new_n3574_ = 1'b1;
default : new_n3574_ = 1'b0;
endcase
casez ({u[2], new_n151_})
2'b01 : new_n3575_ = 1'b1;
default : new_n3575_ = 1'b0;
endcase
casez ({new_n97_, new_n152_})
2'b11 : new_n3576_ = 1'b1;
default : new_n3576_ = 1'b0;
endcase
casez ({new_n103_, new_n153_})
2'b11 : new_n3577_ = 1'b1;
default : new_n3577_ = 1'b0;
endcase
casez ({u[2], new_n158_})
2'b11 : new_n3578_ = 1'b1;
default : new_n3578_ = 1'b0;
endcase
casez ({new_n80_, new_n158_})
2'b11 : new_n3579_ = 1'b1;
default : new_n3579_ = 1'b0;
endcase
casez ({new_n80_, new_n159_})
2'b11 : new_n3580_ = 1'b1;
default : new_n3580_ = 1'b0;
endcase
casez ({new_n85_, new_n162_})
2'b11 : new_n3581_ = 1'b1;
default : new_n3581_ = 1'b0;
endcase
casez ({new_n98_, new_n163_})
2'b11 : new_n3582_ = 1'b1;
default : new_n3582_ = 1'b0;
endcase
casez ({new_n92_, new_n167_})
2'b11 : new_n3583_ = 1'b1;
default : new_n3583_ = 1'b0;
endcase
casez ({new_n80_, new_n167_})
2'b11 : new_n3584_ = 1'b1;
default : new_n3584_ = 1'b0;
endcase
casez ({new_n93_, new_n167_})
2'b11 : new_n3585_ = 1'b1;
default : new_n3585_ = 1'b0;
endcase
casez ({new_n79_, new_n174_})
2'b11 : new_n3586_ = 1'b1;
default : new_n3586_ = 1'b0;
endcase
casez ({new_n80_, new_n177_})
2'b11 : new_n3587_ = 1'b1;
default : new_n3587_ = 1'b0;
endcase
casez ({new_n92_, new_n178_})
2'b11 : new_n3588_ = 1'b1;
default : new_n3588_ = 1'b0;
endcase
casez ({new_n80_, new_n180_})
2'b11 : new_n3589_ = 1'b1;
default : new_n3589_ = 1'b0;
endcase
casez ({new_n92_, new_n199_})
2'b11 : new_n3590_ = 1'b1;
default : new_n3590_ = 1'b0;
endcase
casez ({new_n97_, new_n205_})
2'b11 : new_n3591_ = 1'b1;
default : new_n3591_ = 1'b0;
endcase
casez ({new_n97_, new_n213_})
2'b11 : new_n3592_ = 1'b1;
default : new_n3592_ = 1'b0;
endcase
casez ({new_n83_, new_n217_})
2'b11 : new_n3593_ = 1'b1;
default : new_n3593_ = 1'b0;
endcase
casez ({new_n84_, new_n218_})
2'b11 : new_n3594_ = 1'b1;
default : new_n3594_ = 1'b0;
endcase
casez ({new_n89_, new_n115_})
2'b11 : new_n3595_ = 1'b1;
default : new_n3595_ = 1'b0;
endcase
casez ({v[2], new_n115_})
2'b11 : new_n3596_ = 1'b1;
default : new_n3596_ = 1'b0;
endcase
casez ({new_n104_, new_n115_})
2'b11 : new_n3597_ = 1'b1;
default : new_n3597_ = 1'b0;
endcase
casez ({new_n88_, new_n116_})
2'b11 : new_n3598_ = 1'b1;
default : new_n3598_ = 1'b0;
endcase
casez ({new_n94_, new_n118_})
2'b11 : new_n3599_ = 1'b1;
default : new_n3599_ = 1'b0;
endcase
casez ({new_n97_, new_n126_})
2'b11 : new_n3600_ = 1'b1;
default : new_n3600_ = 1'b0;
endcase
casez ({u[2], new_n128_})
2'b11 : new_n3601_ = 1'b1;
default : new_n3601_ = 1'b0;
endcase
casez ({v[0], new_n131_})
2'b01 : new_n3602_ = 1'b1;
default : new_n3602_ = 1'b0;
endcase
casez ({new_n210_, new_n754_, new_n397_, new_n3602_})
4'b11?? : new_n3603_ = 1'b1;
4'b??11 : new_n3603_ = 1'b1;
default : new_n3603_ = 1'b0;
endcase
casez ({new_n104_, new_n130_})
2'b11 : new_n3604_ = 1'b1;
default : new_n3604_ = 1'b0;
endcase
casez ({new_n89_, new_n133_})
2'b11 : new_n3605_ = 1'b1;
default : new_n3605_ = 1'b0;
endcase
casez ({new_n83_, new_n137_})
2'b11 : new_n3606_ = 1'b1;
default : new_n3606_ = 1'b0;
endcase
casez ({new_n88_, new_n139_})
2'b11 : new_n3607_ = 1'b1;
default : new_n3607_ = 1'b0;
endcase
casez ({new_n95_, new_n139_})
2'b11 : new_n3608_ = 1'b1;
default : new_n3608_ = 1'b0;
endcase
casez ({x[2], new_n139_})
2'b11 : new_n3609_ = 1'b1;
default : new_n3609_ = 1'b0;
endcase
casez ({new_n126_, new_n265_})
2'b00 : new_n3610_ = 1'b1;
default : new_n3610_ = 1'b0;
endcase
casez ({new_n89_, new_n295_, new_n1901_})
3'b01? : new_n3611_ = 1'b1;
3'b??1 : new_n3611_ = 1'b1;
default : new_n3611_ = 1'b0;
endcase
casez ({new_n92_, new_n763_, new_n350_})
3'b11? : new_n3612_ = 1'b1;
3'b??1 : new_n3612_ = 1'b1;
default : new_n3612_ = 1'b0;
endcase
casez ({new_n219_, new_n763_, new_n223_, new_n604_})
4'b11?? : new_n3613_ = 1'b1;
4'b??11 : new_n3613_ = 1'b1;
default : new_n3613_ = 1'b0;
endcase
casez ({new_n244_, new_n480_})
2'b00 : new_n3614_ = 1'b1;
default : new_n3614_ = 1'b0;
endcase
casez ({new_n115_, new_n341_, new_n430_, new_n764_})
4'b11?? : new_n3615_ = 1'b1;
4'b??11 : new_n3615_ = 1'b1;
default : new_n3615_ = 1'b0;
endcase
casez ({new_n710_, new_n1143_})
2'b00 : new_n3616_ = 1'b1;
default : new_n3616_ = 1'b0;
endcase
casez ({new_n96_, new_n261_, new_n481_})
3'b01? : new_n3617_ = 1'b1;
3'b??1 : new_n3617_ = 1'b1;
default : new_n3617_ = 1'b0;
endcase
casez ({new_n4633_, new_n1903_})
2'b1? : new_n3618_ = 1'b1;
2'b?1 : new_n3618_ = 1'b1;
default : new_n3618_ = 1'b0;
endcase
casez ({new_n153_, new_n166_, new_n1903_})
3'b11? : new_n3619_ = 1'b1;
3'b??1 : new_n3619_ = 1'b1;
default : new_n3619_ = 1'b0;
endcase
casez ({v[1], new_n265_, new_n1904_})
3'b01? : new_n3620_ = 1'b1;
3'b??1 : new_n3620_ = 1'b1;
default : new_n3620_ = 1'b0;
endcase
casez ({new_n1142_, new_n1144_})
2'b00 : new_n3621_ = 1'b1;
default : new_n3621_ = 1'b0;
endcase
casez ({new_n378_, new_n481_})
2'b00 : new_n3622_ = 1'b1;
default : new_n3622_ = 1'b0;
endcase
casez ({x[0], new_n103_, new_n275_, new_n1906_})
4'b001? : new_n3623_ = 1'b1;
4'b???1 : new_n3623_ = 1'b1;
default : new_n3623_ = 1'b0;
endcase
casez ({new_n1118_, new_n1906_})
2'b00 : new_n3624_ = 1'b1;
default : new_n3624_ = 1'b0;
endcase
casez ({new_n96_, new_n122_, new_n768_})
3'b11? : new_n3625_ = 1'b1;
3'b??1 : new_n3625_ = 1'b1;
default : new_n3625_ = 1'b0;
endcase
casez ({new_n1856_, new_n1908_})
2'b00 : new_n3626_ = 1'b1;
default : new_n3626_ = 1'b0;
endcase
casez ({y[2], new_n236_, new_n1147_})
3'b11? : new_n3627_ = 1'b1;
3'b??1 : new_n3627_ = 1'b1;
default : new_n3627_ = 1'b0;
endcase
casez ({new_n538_, new_n1145_})
2'b00 : new_n3628_ = 1'b1;
default : new_n3628_ = 1'b0;
endcase
casez ({new_n1895_, new_n1908_})
2'b00 : new_n3629_ = 1'b1;
default : new_n3629_ = 1'b0;
endcase
casez ({new_n602_, new_n1909_})
2'b00 : new_n3630_ = 1'b1;
default : new_n3630_ = 1'b0;
endcase
casez ({new_n336_, new_n1909_})
2'b00 : new_n3631_ = 1'b1;
default : new_n3631_ = 1'b0;
endcase
casez ({new_n4633_, new_n1910_})
2'b1? : new_n3632_ = 1'b1;
2'b?1 : new_n3632_ = 1'b1;
default : new_n3632_ = 1'b0;
endcase
casez ({new_n259_, new_n1146_})
2'b00 : new_n3633_ = 1'b1;
default : new_n3633_ = 1'b0;
endcase
casez ({new_n956_, new_n1911_})
2'b00 : new_n3634_ = 1'b1;
default : new_n3634_ = 1'b0;
endcase
casez ({new_n214_, new_n320_, new_n482_})
3'b10? : new_n3635_ = 1'b1;
3'b??1 : new_n3635_ = 1'b1;
default : new_n3635_ = 1'b0;
endcase
casez ({new_n1339_, new_n1912_})
2'b00 : new_n3636_ = 1'b1;
default : new_n3636_ = 1'b0;
endcase
casez ({u[1], new_n482_, new_n4649_})
3'b01? : new_n3637_ = 1'b1;
3'b??1 : new_n3637_ = 1'b1;
default : new_n3637_ = 1'b0;
endcase
casez ({new_n740_, new_n1913_})
2'b00 : new_n3638_ = 1'b1;
default : new_n3638_ = 1'b0;
endcase
casez ({new_n718_, new_n1916_})
2'b00 : new_n3639_ = 1'b1;
default : new_n3639_ = 1'b0;
endcase
casez ({new_n160_, new_n615_, new_n1149_})
3'b10? : new_n3640_ = 1'b1;
3'b??1 : new_n3640_ = 1'b1;
default : new_n3640_ = 1'b0;
endcase
casez ({new_n797_, new_n1917_})
2'b00 : new_n3641_ = 1'b1;
default : new_n3641_ = 1'b0;
endcase
casez ({new_n1891_, new_n1917_})
2'b00 : new_n3642_ = 1'b1;
default : new_n3642_ = 1'b0;
endcase
casez ({new_n196_, new_n774_})
2'b01 : new_n3643_ = 1'b1;
default : new_n3643_ = 1'b0;
endcase
casez ({new_n1017_, new_n1918_})
2'b00 : new_n3644_ = 1'b1;
default : new_n3644_ = 1'b0;
endcase
casez ({new_n191_, new_n764_, new_n1150_})
3'b11? : new_n3645_ = 1'b1;
3'b??1 : new_n3645_ = 1'b1;
default : new_n3645_ = 1'b0;
endcase
casez ({new_n540_, new_n1921_})
2'b00 : new_n3646_ = 1'b1;
default : new_n3646_ = 1'b0;
endcase
casez ({new_n619_, new_n1263_, new_n1923_})
3'b10? : new_n3647_ = 1'b1;
3'b??1 : new_n3647_ = 1'b1;
default : new_n3647_ = 1'b0;
endcase
casez ({new_n789_, new_n1923_})
2'b00 : new_n3648_ = 1'b1;
default : new_n3648_ = 1'b0;
endcase
casez ({new_n1374_, new_n1923_})
2'b00 : new_n3649_ = 1'b1;
default : new_n3649_ = 1'b0;
endcase
casez ({new_n107_, new_n405_, new_n1924_})
3'b01? : new_n3650_ = 1'b1;
3'b??1 : new_n3650_ = 1'b1;
default : new_n3650_ = 1'b0;
endcase
casez ({u[1], new_n776_, new_n377_})
3'b11? : new_n3651_ = 1'b1;
3'b0?1 : new_n3651_ = 1'b1;
default : new_n3651_ = 1'b0;
endcase
casez ({u[1], new_n372_, new_n265_, new_n487_})
4'b01?? : new_n3652_ = 1'b1;
4'b??11 : new_n3652_ = 1'b1;
default : new_n3652_ = 1'b0;
endcase
casez ({new_n1158_, new_n1925_})
2'b00 : new_n3653_ = 1'b1;
default : new_n3653_ = 1'b0;
endcase
casez ({y[2], new_n127_, new_n1925_})
3'b01? : new_n3654_ = 1'b1;
3'b??1 : new_n3654_ = 1'b1;
default : new_n3654_ = 1'b0;
endcase
casez ({new_n154_, new_n258_, new_n777_})
3'b11? : new_n3655_ = 1'b1;
3'b??1 : new_n3655_ = 1'b1;
default : new_n3655_ = 1'b0;
endcase
casez ({new_n4658_, new_n215_, new_n487_})
3'b1?? : new_n3656_ = 1'b1;
3'b?11 : new_n3656_ = 1'b1;
default : new_n3656_ = 1'b0;
endcase
casez ({new_n214_, new_n229_, new_n1152_})
3'b11? : new_n3657_ = 1'b1;
3'b??1 : new_n3657_ = 1'b1;
default : new_n3657_ = 1'b0;
endcase
casez ({new_n118_, new_n228_, new_n1927_})
3'b11? : new_n3658_ = 1'b1;
3'b??1 : new_n3658_ = 1'b1;
default : new_n3658_ = 1'b0;
endcase
casez ({new_n86_, new_n222_, new_n1153_})
3'b11? : new_n3659_ = 1'b1;
3'b??1 : new_n3659_ = 1'b1;
default : new_n3659_ = 1'b0;
endcase
casez ({new_n937_, new_n1153_})
2'b00 : new_n3660_ = 1'b1;
default : new_n3660_ = 1'b0;
endcase
casez ({new_n90_, new_n194_, new_n175_, new_n489_})
4'b11?? : new_n3661_ = 1'b1;
4'b??11 : new_n3661_ = 1'b1;
default : new_n3661_ = 1'b0;
endcase
casez ({new_n204_, new_n249_, new_n1930_})
3'b11? : new_n3662_ = 1'b1;
3'b??1 : new_n3662_ = 1'b1;
default : new_n3662_ = 1'b0;
endcase
casez ({new_n1875_, new_n1930_})
2'b00 : new_n3663_ = 1'b1;
default : new_n3663_ = 1'b0;
endcase
casez ({y[2], new_n205_, new_n1932_})
3'b11? : new_n3664_ = 1'b1;
3'b??1 : new_n3664_ = 1'b1;
default : new_n3664_ = 1'b0;
endcase
casez ({new_n301_, new_n478_, new_n1154_})
3'b11? : new_n3665_ = 1'b1;
3'b??1 : new_n3665_ = 1'b1;
default : new_n3665_ = 1'b0;
endcase
casez ({new_n361_, new_n1932_})
2'b00 : new_n3666_ = 1'b1;
default : new_n3666_ = 1'b0;
endcase
casez ({new_n1560_, new_n1933_})
2'b00 : new_n3667_ = 1'b1;
default : new_n3667_ = 1'b0;
endcase
casez ({new_n220_, new_n491_})
2'b01 : new_n3668_ = 1'b1;
default : new_n3668_ = 1'b0;
endcase
casez ({new_n134_, new_n398_, new_n778_})
3'b11? : new_n3669_ = 1'b1;
3'b??1 : new_n3669_ = 1'b1;
default : new_n3669_ = 1'b0;
endcase
casez ({new_n1130_, new_n1933_})
2'b00 : new_n3670_ = 1'b1;
default : new_n3670_ = 1'b0;
endcase
casez ({new_n198_, new_n493_})
2'b00 : new_n3671_ = 1'b1;
default : new_n3671_ = 1'b0;
endcase
casez ({u[1], new_n388_, new_n85_, new_n493_})
4'b01?? : new_n3672_ = 1'b1;
4'b??11 : new_n3672_ = 1'b1;
default : new_n3672_ = 1'b0;
endcase
casez ({new_n274_, new_n493_})
2'b00 : new_n3673_ = 1'b1;
default : new_n3673_ = 1'b0;
endcase
casez ({new_n91_, new_n118_, new_n279_, new_n493_})
4'b11?? : new_n3674_ = 1'b1;
4'b??11 : new_n3674_ = 1'b1;
default : new_n3674_ = 1'b0;
endcase
casez ({new_n101_, new_n1935_, new_n1596_})
3'b11? : new_n3675_ = 1'b1;
3'b??1 : new_n3675_ = 1'b1;
default : new_n3675_ = 1'b0;
endcase
casez ({new_n207_, new_n493_})
2'b00 : new_n3676_ = 1'b1;
default : new_n3676_ = 1'b0;
endcase
casez ({new_n293_, new_n444_, new_n779_})
3'b11? : new_n3677_ = 1'b1;
3'b??1 : new_n3677_ = 1'b1;
default : new_n3677_ = 1'b0;
endcase
casez ({new_n221_, new_n224_, new_n1936_})
3'b11? : new_n3678_ = 1'b1;
3'b??1 : new_n3678_ = 1'b1;
default : new_n3678_ = 1'b0;
endcase
casez ({new_n145_, new_n429_, new_n360_, new_n494_})
4'b11?? : new_n3679_ = 1'b1;
4'b??11 : new_n3679_ = 1'b1;
default : new_n3679_ = 1'b0;
endcase
casez ({new_n678_, new_n1936_})
2'b00 : new_n3680_ = 1'b1;
default : new_n3680_ = 1'b0;
endcase
casez ({new_n868_, new_n1156_})
2'b00 : new_n3681_ = 1'b1;
default : new_n3681_ = 1'b0;
endcase
casez ({new_n208_, new_n364_, new_n1936_})
3'b10? : new_n3682_ = 1'b1;
3'b??1 : new_n3682_ = 1'b1;
default : new_n3682_ = 1'b0;
endcase
casez ({new_n94_, new_n494_, new_n122_, new_n407_})
4'b11?? : new_n3683_ = 1'b1;
4'b??11 : new_n3683_ = 1'b1;
default : new_n3683_ = 1'b0;
endcase
casez ({new_n88_, new_n366_, new_n779_})
3'b01? : new_n3684_ = 1'b1;
3'b??1 : new_n3684_ = 1'b1;
default : new_n3684_ = 1'b0;
endcase
casez ({new_n247_, new_n441_, new_n320_, new_n494_})
4'b11?? : new_n3685_ = 1'b1;
4'b??01 : new_n3685_ = 1'b1;
default : new_n3685_ = 1'b0;
endcase
casez ({new_n85_, new_n287_, new_n1939_})
3'b11? : new_n3686_ = 1'b1;
3'b??1 : new_n3686_ = 1'b1;
default : new_n3686_ = 1'b0;
endcase
casez ({new_n951_, new_n1157_})
2'b00 : new_n3687_ = 1'b1;
default : new_n3687_ = 1'b0;
endcase
casez ({new_n502_, new_n1940_})
2'b00 : new_n3688_ = 1'b1;
default : new_n3688_ = 1'b0;
endcase
casez ({new_n222_, new_n495_})
2'b00 : new_n3689_ = 1'b1;
default : new_n3689_ = 1'b0;
endcase
casez ({new_n190_, new_n1941_})
2'b00 : new_n3690_ = 1'b1;
default : new_n3690_ = 1'b0;
endcase
casez ({new_n742_, new_n1942_})
2'b00 : new_n3691_ = 1'b1;
default : new_n3691_ = 1'b0;
endcase
casez ({new_n97_, new_n496_, new_n177_, new_n309_})
4'b11?? : new_n3692_ = 1'b1;
4'b??11 : new_n3692_ = 1'b1;
default : new_n3692_ = 1'b0;
endcase
casez ({new_n1370_, new_n1943_})
2'b00 : new_n3693_ = 1'b1;
default : new_n3693_ = 1'b0;
endcase
casez ({new_n717_, new_n1158_})
2'b00 : new_n3694_ = 1'b1;
default : new_n3694_ = 1'b0;
endcase
casez ({new_n778_, new_n780_})
2'b00 : new_n3695_ = 1'b1;
default : new_n3695_ = 1'b0;
endcase
casez ({new_n4585_, new_n382_})
2'b1? : new_n3696_ = 1'b1;
2'b?1 : new_n3696_ = 1'b1;
default : new_n3696_ = 1'b0;
endcase
casez ({new_n4583_, new_n166_, new_n719_})
3'b1?? : new_n3697_ = 1'b1;
3'b?11 : new_n3697_ = 1'b1;
default : new_n3697_ = 1'b0;
endcase
casez ({new_n768_, new_n1159_})
2'b00 : new_n3698_ = 1'b1;
default : new_n3698_ = 1'b0;
endcase
casez ({new_n280_, new_n1945_})
2'b00 : new_n3699_ = 1'b1;
default : new_n3699_ = 1'b0;
endcase
casez ({new_n673_, new_n1945_})
2'b00 : new_n3700_ = 1'b1;
default : new_n3700_ = 1'b0;
endcase
casez ({new_n1885_, new_n1946_})
2'b00 : new_n3701_ = 1'b1;
default : new_n3701_ = 1'b0;
endcase
casez ({new_n83_, new_n116_, new_n1947_})
3'b01? : new_n3702_ = 1'b1;
3'b??1 : new_n3702_ = 1'b1;
default : new_n3702_ = 1'b0;
endcase
casez ({new_n863_, new_n1947_})
2'b00 : new_n3703_ = 1'b1;
default : new_n3703_ = 1'b0;
endcase
casez ({new_n144_, new_n749_, new_n235_, new_n1160_})
4'b11?? : new_n3704_ = 1'b1;
4'b??11 : new_n3704_ = 1'b1;
default : new_n3704_ = 1'b0;
endcase
casez ({new_n199_, new_n497_})
2'b00 : new_n3705_ = 1'b1;
default : new_n3705_ = 1'b0;
endcase
casez ({new_n1172_, new_n1948_})
2'b00 : new_n3706_ = 1'b1;
default : new_n3706_ = 1'b0;
endcase
casez ({v[1], new_n1949_, new_n1010_})
3'b11? : new_n3707_ = 1'b1;
3'b??1 : new_n3707_ = 1'b1;
default : new_n3707_ = 1'b0;
endcase
casez ({new_n1162_, new_n1949_})
2'b00 : new_n3708_ = 1'b1;
default : new_n3708_ = 1'b0;
endcase
casez ({new_n792_, new_n1950_})
2'b00 : new_n3709_ = 1'b1;
default : new_n3709_ = 1'b0;
endcase
casez ({x[0], new_n1950_, new_n97_, new_n1386_})
4'b01?? : new_n3710_ = 1'b1;
4'b??11 : new_n3710_ = 1'b1;
default : new_n3710_ = 1'b0;
endcase
casez ({new_n268_, new_n1951_})
2'b00 : new_n3711_ = 1'b1;
default : new_n3711_ = 1'b0;
endcase
casez ({y[1], new_n783_, v[2], new_n430_})
4'b01?? : new_n3712_ = 1'b1;
4'b??01 : new_n3712_ = 1'b1;
default : new_n3712_ = 1'b0;
endcase
casez ({new_n109_, new_n397_, new_n498_})
3'b01? : new_n3713_ = 1'b1;
3'b??1 : new_n3713_ = 1'b1;
default : new_n3713_ = 1'b0;
endcase
casez ({x[2], new_n398_, new_n1952_})
3'b01? : new_n3714_ = 1'b1;
3'b??1 : new_n3714_ = 1'b1;
default : new_n3714_ = 1'b0;
endcase
casez ({new_n86_, new_n381_, new_n1953_})
3'b11? : new_n3715_ = 1'b1;
3'b??1 : new_n3715_ = 1'b1;
default : new_n3715_ = 1'b0;
endcase
casez ({new_n454_, new_n498_})
2'b00 : new_n3716_ = 1'b1;
default : new_n3716_ = 1'b0;
endcase
casez ({new_n792_, new_n1954_})
2'b00 : new_n3717_ = 1'b1;
default : new_n3717_ = 1'b0;
endcase
casez ({x[2], new_n1955_, new_n1630_})
3'b01? : new_n3718_ = 1'b1;
3'b??1 : new_n3718_ = 1'b1;
default : new_n3718_ = 1'b0;
endcase
casez ({new_n497_, new_n498_})
2'b00 : new_n3719_ = 1'b1;
default : new_n3719_ = 1'b0;
endcase
casez ({new_n356_, new_n1955_})
2'b00 : new_n3720_ = 1'b1;
default : new_n3720_ = 1'b0;
endcase
casez ({new_n1630_, new_n1956_})
2'b00 : new_n3721_ = 1'b1;
default : new_n3721_ = 1'b0;
endcase
casez ({new_n89_, new_n310_, new_n1164_})
3'b11? : new_n3722_ = 1'b1;
3'b??1 : new_n3722_ = 1'b1;
default : new_n3722_ = 1'b0;
endcase
casez ({new_n1388_, new_n1956_})
2'b00 : new_n3723_ = 1'b1;
default : new_n3723_ = 1'b0;
endcase
casez ({new_n211_, new_n346_, new_n498_})
3'b11? : new_n3724_ = 1'b1;
3'b??1 : new_n3724_ = 1'b1;
default : new_n3724_ = 1'b0;
endcase
casez ({new_n636_, new_n1165_})
2'b00 : new_n3725_ = 1'b1;
default : new_n3725_ = 1'b0;
endcase
casez ({new_n946_, new_n1164_})
2'b00 : new_n3726_ = 1'b1;
default : new_n3726_ = 1'b0;
endcase
casez ({new_n83_, new_n499_, new_n405_})
3'b11? : new_n3727_ = 1'b1;
3'b??1 : new_n3727_ = 1'b1;
default : new_n3727_ = 1'b0;
endcase
casez ({new_n182_, new_n319_, new_n215_, new_n499_})
4'b10?? : new_n3728_ = 1'b1;
4'b??11 : new_n3728_ = 1'b1;
default : new_n3728_ = 1'b0;
endcase
casez ({new_n767_, new_n1164_})
2'b00 : new_n3729_ = 1'b1;
default : new_n3729_ = 1'b0;
endcase
casez ({new_n118_, new_n196_, new_n785_})
3'b11? : new_n3730_ = 1'b1;
3'b??1 : new_n3730_ = 1'b1;
default : new_n3730_ = 1'b0;
endcase
casez ({new_n779_, new_n785_})
2'b00 : new_n3731_ = 1'b1;
default : new_n3731_ = 1'b0;
endcase
casez ({new_n89_, new_n1165_, new_n221_, new_n599_})
4'b01?? : new_n3732_ = 1'b1;
4'b??11 : new_n3732_ = 1'b1;
default : new_n3732_ = 1'b0;
endcase
casez ({new_n448_, new_n1958_})
2'b00 : new_n3733_ = 1'b1;
default : new_n3733_ = 1'b0;
endcase
casez ({new_n4590_, new_n785_})
2'b1? : new_n3734_ = 1'b1;
2'b?1 : new_n3734_ = 1'b1;
default : new_n3734_ = 1'b0;
endcase
casez ({new_n742_, new_n1961_})
2'b00 : new_n3735_ = 1'b1;
default : new_n3735_ = 1'b0;
endcase
casez ({new_n265_, new_n501_})
2'b00 : new_n3736_ = 1'b1;
default : new_n3736_ = 1'b0;
endcase
casez ({u[1], new_n541_, new_n1961_})
3'b01? : new_n3737_ = 1'b1;
3'b??1 : new_n3737_ = 1'b1;
default : new_n3737_ = 1'b0;
endcase
casez ({new_n497_, new_n501_})
2'b00 : new_n3738_ = 1'b1;
default : new_n3738_ = 1'b0;
endcase
casez ({new_n873_, new_n1962_})
2'b00 : new_n3739_ = 1'b1;
default : new_n3739_ = 1'b0;
endcase
casez ({new_n131_, new_n629_, new_n616_, new_n786_})
4'b10?? : new_n3740_ = 1'b1;
4'b??11 : new_n3740_ = 1'b1;
default : new_n3740_ = 1'b0;
endcase
casez ({new_n109_, new_n787_, new_n154_, new_n222_})
4'b01?? : new_n3741_ = 1'b1;
4'b??11 : new_n3741_ = 1'b1;
default : new_n3741_ = 1'b0;
endcase
casez ({y[2], new_n121_, new_n787_})
3'b11? : new_n3742_ = 1'b1;
3'b??1 : new_n3742_ = 1'b1;
default : new_n3742_ = 1'b0;
endcase
casez ({u[0], new_n669_, new_n83_, new_n1168_})
4'b01?? : new_n3743_ = 1'b1;
4'b??01 : new_n3743_ = 1'b1;
default : new_n3743_ = 1'b0;
endcase
casez ({new_n104_, new_n489_, new_n1963_})
3'b11? : new_n3744_ = 1'b1;
3'b??1 : new_n3744_ = 1'b1;
default : new_n3744_ = 1'b0;
endcase
casez ({new_n93_, new_n281_, new_n501_})
3'b01? : new_n3745_ = 1'b1;
3'b??1 : new_n3745_ = 1'b1;
default : new_n3745_ = 1'b0;
endcase
casez ({new_n423_, new_n1964_})
2'b00 : new_n3746_ = 1'b1;
default : new_n3746_ = 1'b0;
endcase
casez ({v[1], new_n205_, new_n787_})
3'b11? : new_n3747_ = 1'b1;
3'b??1 : new_n3747_ = 1'b1;
default : new_n3747_ = 1'b0;
endcase
casez ({new_n550_, new_n1168_})
2'b10 : new_n3748_ = 1'b1;
default : new_n3748_ = 1'b0;
endcase
casez ({new_n144_, new_n502_})
2'b00 : new_n3749_ = 1'b1;
default : new_n3749_ = 1'b0;
endcase
casez ({new_n295_, new_n788_})
2'b00 : new_n3750_ = 1'b1;
default : new_n3750_ = 1'b0;
endcase
casez ({new_n289_, new_n1169_})
2'b00 : new_n3751_ = 1'b1;
default : new_n3751_ = 1'b0;
endcase
casez ({new_n84_, new_n511_, new_n1170_})
3'b10? : new_n3752_ = 1'b1;
3'b??1 : new_n3752_ = 1'b1;
default : new_n3752_ = 1'b0;
endcase
casez ({new_n185_, new_n503_})
2'b00 : new_n3753_ = 1'b1;
default : new_n3753_ = 1'b0;
endcase
casez ({new_n87_, new_n294_, new_n445_, new_n503_})
4'b11?? : new_n3754_ = 1'b1;
4'b??11 : new_n3754_ = 1'b1;
default : new_n3754_ = 1'b0;
endcase
casez ({new_n496_, new_n503_})
2'b00 : new_n3755_ = 1'b1;
default : new_n3755_ = 1'b0;
endcase
casez ({new_n97_, new_n244_, new_n1170_})
3'b11? : new_n3756_ = 1'b1;
3'b??1 : new_n3756_ = 1'b1;
default : new_n3756_ = 1'b0;
endcase
casez ({new_n94_, new_n961_, new_n428_, new_n1171_})
4'b11?? : new_n3757_ = 1'b1;
4'b??01 : new_n3757_ = 1'b1;
default : new_n3757_ = 1'b0;
endcase
casez ({new_n154_, new_n271_, new_n481_, new_n1171_})
4'b11?? : new_n3758_ = 1'b1;
4'b??11 : new_n3758_ = 1'b1;
default : new_n3758_ = 1'b0;
endcase
casez ({new_n671_, new_n1172_})
2'b00 : new_n3759_ = 1'b1;
default : new_n3759_ = 1'b0;
endcase
casez ({new_n600_, new_n789_})
2'b00 : new_n3760_ = 1'b1;
default : new_n3760_ = 1'b0;
endcase
casez ({new_n782_, new_n789_})
2'b00 : new_n3761_ = 1'b1;
default : new_n3761_ = 1'b0;
endcase
casez ({new_n4587_, new_n148_, new_n542_})
3'b1?? : new_n3762_ = 1'b1;
3'b?11 : new_n3762_ = 1'b1;
default : new_n3762_ = 1'b0;
endcase
casez ({new_n85_, new_n619_, new_n1175_})
3'b11? : new_n3763_ = 1'b1;
3'b??1 : new_n3763_ = 1'b1;
default : new_n3763_ = 1'b0;
endcase
casez ({new_n1135_, new_n1176_})
2'b00 : new_n3764_ = 1'b1;
default : new_n3764_ = 1'b0;
endcase
casez ({new_n83_, new_n240_, new_n792_})
3'b11? : new_n3765_ = 1'b1;
3'b??1 : new_n3765_ = 1'b1;
default : new_n3765_ = 1'b0;
endcase
casez ({new_n743_, new_n1176_})
2'b00 : new_n3766_ = 1'b1;
default : new_n3766_ = 1'b0;
endcase
casez ({new_n496_, new_n1177_})
2'b00 : new_n3767_ = 1'b1;
default : new_n3767_ = 1'b0;
endcase
casez ({new_n424_, new_n793_})
2'b00 : new_n3768_ = 1'b1;
default : new_n3768_ = 1'b0;
endcase
casez ({x[0], new_n952_, new_n1178_})
3'b11? : new_n3769_ = 1'b1;
3'b??1 : new_n3769_ = 1'b1;
default : new_n3769_ = 1'b0;
endcase
casez ({new_n205_, new_n1179_, new_n267_, new_n282_})
4'b11?? : new_n3770_ = 1'b1;
4'b??11 : new_n3770_ = 1'b1;
default : new_n3770_ = 1'b0;
endcase
casez ({new_n538_, new_n793_})
2'b00 : new_n3771_ = 1'b1;
default : new_n3771_ = 1'b0;
endcase
casez ({new_n383_, new_n1180_})
2'b00 : new_n3772_ = 1'b1;
default : new_n3772_ = 1'b0;
endcase
casez ({new_n407_, new_n1180_})
2'b00 : new_n3773_ = 1'b1;
default : new_n3773_ = 1'b0;
endcase
casez ({new_n4669_, new_n189_, new_n264_})
3'b1?? : new_n3774_ = 1'b1;
3'b?11 : new_n3774_ = 1'b1;
default : new_n3774_ = 1'b0;
endcase
casez ({new_n323_, new_n793_})
2'b00 : new_n3775_ = 1'b1;
default : new_n3775_ = 1'b0;
endcase
casez ({new_n718_, new_n1180_})
2'b00 : new_n3776_ = 1'b1;
default : new_n3776_ = 1'b0;
endcase
casez ({new_n104_, new_n398_, new_n1180_})
3'b11? : new_n3777_ = 1'b1;
3'b??1 : new_n3777_ = 1'b1;
default : new_n3777_ = 1'b0;
endcase
casez ({new_n86_, new_n388_, new_n1181_})
3'b11? : new_n3778_ = 1'b1;
3'b??1 : new_n3778_ = 1'b1;
default : new_n3778_ = 1'b0;
endcase
casez ({new_n1180_, new_n1181_})
2'b00 : new_n3779_ = 1'b1;
default : new_n3779_ = 1'b0;
endcase
casez ({new_n183_, new_n212_, new_n238_, new_n796_})
4'b11?? : new_n3780_ = 1'b1;
4'b??11 : new_n3780_ = 1'b1;
default : new_n3780_ = 1'b0;
endcase
casez ({new_n524_, new_n796_, new_n619_, new_n744_})
4'b11?? : new_n3781_ = 1'b1;
4'b??11 : new_n3781_ = 1'b1;
default : new_n3781_ = 1'b0;
endcase
casez ({new_n350_, new_n797_})
2'b00 : new_n3782_ = 1'b1;
default : new_n3782_ = 1'b0;
endcase
casez ({new_n152_, new_n265_})
2'b00 : new_n3783_ = 1'b1;
default : new_n3783_ = 1'b0;
endcase
casez ({new_n261_, new_n799_, new_n302_, new_n391_})
4'b11?? : new_n3784_ = 1'b1;
4'b??01 : new_n3784_ = 1'b1;
default : new_n3784_ = 1'b0;
endcase
casez ({x[1], new_n799_, new_n718_})
3'b01? : new_n3785_ = 1'b1;
3'b??1 : new_n3785_ = 1'b1;
default : new_n3785_ = 1'b0;
endcase
casez ({new_n96_, new_n267_, new_n217_})
3'b01? : new_n3786_ = 1'b1;
3'b??1 : new_n3786_ = 1'b1;
default : new_n3786_ = 1'b0;
endcase
casez ({new_n183_, new_n523_})
2'b01 : new_n3787_ = 1'b1;
default : new_n3787_ = 1'b0;
endcase
casez ({u[1], new_n524_, new_n230_, new_n337_})
4'b11?? : new_n3788_ = 1'b1;
4'b??11 : new_n3788_ = 1'b1;
default : new_n3788_ = 1'b0;
endcase
casez ({new_n424_, new_n525_})
2'b00 : new_n3789_ = 1'b1;
default : new_n3789_ = 1'b0;
endcase
casez ({new_n334_, new_n525_})
2'b00 : new_n3790_ = 1'b1;
default : new_n3790_ = 1'b0;
endcase
casez ({new_n4588_, v[0], new_n408_})
3'b1?? : new_n3791_ = 1'b1;
3'b?11 : new_n3791_ = 1'b1;
default : new_n3791_ = 1'b0;
endcase
casez ({new_n377_, new_n526_})
2'b00 : new_n3792_ = 1'b1;
default : new_n3792_ = 1'b0;
endcase
casez ({new_n88_, new_n131_, new_n527_})
3'b11? : new_n3793_ = 1'b1;
3'b??1 : new_n3793_ = 1'b1;
default : new_n3793_ = 1'b0;
endcase
casez ({new_n4631_, new_n369_, new_n530_})
3'b1?? : new_n3794_ = 1'b1;
3'b?11 : new_n3794_ = 1'b1;
default : new_n3794_ = 1'b0;
endcase
casez ({new_n145_, new_n237_, new_n181_, new_n271_})
4'b11?? : new_n3795_ = 1'b1;
4'b??01 : new_n3795_ = 1'b1;
default : new_n3795_ = 1'b0;
endcase
casez ({v[2], new_n96_, new_n271_})
3'b01? : new_n3796_ = 1'b1;
3'b??1 : new_n3796_ = 1'b1;
default : new_n3796_ = 1'b0;
endcase
casez ({new_n190_, new_n417_, new_n535_})
3'b11? : new_n3797_ = 1'b1;
3'b??1 : new_n3797_ = 1'b1;
default : new_n3797_ = 1'b0;
endcase
casez ({new_n360_, new_n488_, new_n535_})
3'b11? : new_n3798_ = 1'b1;
3'b??1 : new_n3798_ = 1'b1;
default : new_n3798_ = 1'b0;
endcase
casez ({new_n4589_, new_n261_, new_n347_})
3'b1?? : new_n3799_ = 1'b1;
3'b?11 : new_n3799_ = 1'b1;
default : new_n3799_ = 1'b0;
endcase
casez ({new_n387_, new_n537_})
2'b00 : new_n3800_ = 1'b1;
default : new_n3800_ = 1'b0;
endcase
casez ({new_n339_, new_n537_})
2'b00 : new_n3801_ = 1'b1;
default : new_n3801_ = 1'b0;
endcase
casez ({y[2], new_n538_, new_n441_})
3'b01? : new_n3802_ = 1'b1;
3'b??1 : new_n3802_ = 1'b1;
default : new_n3802_ = 1'b0;
endcase
casez ({y[2], new_n538_, new_n455_})
3'b11? : new_n3803_ = 1'b1;
3'b??1 : new_n3803_ = 1'b1;
default : new_n3803_ = 1'b0;
endcase
casez ({new_n120_, new_n539_})
2'b00 : new_n3804_ = 1'b1;
default : new_n3804_ = 1'b0;
endcase
casez ({x[0], new_n137_, u[0], new_n157_})
4'b11?? : new_n3805_ = 1'b1;
4'b??11 : new_n3805_ = 1'b1;
default : new_n3805_ = 1'b0;
endcase
casez ({new_n384_, new_n540_})
2'b00 : new_n3806_ = 1'b1;
default : new_n3806_ = 1'b0;
endcase
casez ({new_n126_, new_n821_, new_n260_, new_n294_})
4'b11?? : new_n3807_ = 1'b1;
4'b??11 : new_n3807_ = 1'b1;
default : new_n3807_ = 1'b0;
endcase
casez ({new_n121_, new_n282_, new_n494_, new_n822_})
4'b11?? : new_n3808_ = 1'b1;
4'b??11 : new_n3808_ = 1'b1;
default : new_n3808_ = 1'b0;
endcase
casez ({new_n101_, new_n382_, new_n540_})
3'b11? : new_n3809_ = 1'b1;
3'b??1 : new_n3809_ = 1'b1;
default : new_n3809_ = 1'b0;
endcase
casez ({new_n123_, new_n541_, new_n154_, new_n240_})
4'b11?? : new_n3810_ = 1'b1;
4'b??11 : new_n3810_ = 1'b1;
default : new_n3810_ = 1'b0;
endcase
casez ({new_n167_, new_n207_, new_n223_, new_n541_})
4'b11?? : new_n3811_ = 1'b1;
4'b??11 : new_n3811_ = 1'b1;
default : new_n3811_ = 1'b0;
endcase
casez ({new_n190_, new_n278_, new_n204_, new_n267_})
4'b11?? : new_n3812_ = 1'b1;
4'b??11 : new_n3812_ = 1'b1;
default : new_n3812_ = 1'b0;
endcase
casez ({new_n98_, new_n549_, new_n456_})
3'b11? : new_n3813_ = 1'b1;
3'b??1 : new_n3813_ = 1'b1;
default : new_n3813_ = 1'b0;
endcase
casez ({new_n240_, new_n358_, new_n854_})
3'b11? : new_n3814_ = 1'b1;
3'b??1 : new_n3814_ = 1'b1;
default : new_n3814_ = 1'b0;
endcase
casez ({new_n79_, new_n278_, new_n855_})
3'b11? : new_n3815_ = 1'b1;
3'b??1 : new_n3815_ = 1'b1;
default : new_n3815_ = 1'b0;
endcase
casez ({new_n86_, new_n92_, new_n855_})
3'b11? : new_n3816_ = 1'b1;
3'b??1 : new_n3816_ = 1'b1;
default : new_n3816_ = 1'b0;
endcase
casez ({new_n182_, new_n855_})
2'b00 : new_n3817_ = 1'b1;
default : new_n3817_ = 1'b0;
endcase
casez ({u[1], new_n389_, new_n856_})
3'b11? : new_n3818_ = 1'b1;
3'b??1 : new_n3818_ = 1'b1;
default : new_n3818_ = 1'b0;
endcase
casez ({new_n127_, new_n211_, new_n553_})
3'b11? : new_n3819_ = 1'b1;
3'b??1 : new_n3819_ = 1'b1;
default : new_n3819_ = 1'b0;
endcase
casez ({new_n79_, new_n196_, new_n554_})
3'b11? : new_n3820_ = 1'b1;
3'b??1 : new_n3820_ = 1'b1;
default : new_n3820_ = 1'b0;
endcase
casez ({new_n424_, new_n554_})
2'b00 : new_n3821_ = 1'b1;
default : new_n3821_ = 1'b0;
endcase
casez ({new_n497_, new_n554_})
2'b00 : new_n3822_ = 1'b1;
default : new_n3822_ = 1'b0;
endcase
casez ({new_n289_, new_n557_})
2'b00 : new_n3823_ = 1'b1;
default : new_n3823_ = 1'b0;
endcase
casez ({new_n212_, new_n235_, new_n860_})
3'b11? : new_n3824_ = 1'b1;
3'b??1 : new_n3824_ = 1'b1;
default : new_n3824_ = 1'b0;
endcase
casez ({new_n788_, new_n859_})
2'b00 : new_n3825_ = 1'b1;
default : new_n3825_ = 1'b0;
endcase
casez ({new_n122_, new_n321_, new_n318_, new_n1257_})
4'b11?? : new_n3826_ = 1'b1;
4'b??11 : new_n3826_ = 1'b1;
default : new_n3826_ = 1'b0;
endcase
casez ({new_n501_, new_n1260_})
2'b00 : new_n3827_ = 1'b1;
default : new_n3827_ = 1'b0;
endcase
casez ({new_n4625_, new_n860_})
2'b1? : new_n3828_ = 1'b1;
2'b?1 : new_n3828_ = 1'b1;
default : new_n3828_ = 1'b0;
endcase
casez ({new_n127_, new_n1264_, new_n1157_})
3'b11? : new_n3829_ = 1'b1;
3'b??1 : new_n3829_ = 1'b1;
default : new_n3829_ = 1'b0;
endcase
casez ({new_n343_, new_n486_, new_n861_})
3'b11? : new_n3830_ = 1'b1;
3'b??1 : new_n3830_ = 1'b1;
default : new_n3830_ = 1'b0;
endcase
casez ({x[0], new_n92_, new_n156_, new_n862_})
4'b101? : new_n3831_ = 1'b1;
4'b???1 : new_n3831_ = 1'b1;
default : new_n3831_ = 1'b0;
endcase
casez ({new_n280_, new_n289_})
2'b00 : new_n3832_ = 1'b1;
default : new_n3832_ = 1'b0;
endcase
casez ({new_n199_, new_n1276_, new_n711_})
3'b10? : new_n3833_ = 1'b1;
3'b??1 : new_n3833_ = 1'b1;
default : new_n3833_ = 1'b0;
endcase
casez ({new_n186_, new_n196_, new_n865_})
3'b11? : new_n3834_ = 1'b1;
3'b??1 : new_n3834_ = 1'b1;
default : new_n3834_ = 1'b0;
endcase
casez ({new_n144_, new_n294_})
2'b00 : new_n3835_ = 1'b1;
default : new_n3835_ = 1'b0;
endcase
casez ({new_n212_, new_n659_, new_n866_})
3'b10? : new_n3836_ = 1'b1;
3'b??1 : new_n3836_ = 1'b1;
default : new_n3836_ = 1'b0;
endcase
casez ({new_n262_, new_n619_, new_n866_})
3'b11? : new_n3837_ = 1'b1;
3'b??1 : new_n3837_ = 1'b1;
default : new_n3837_ = 1'b0;
endcase
casez ({new_n145_, new_n674_, new_n867_})
3'b11? : new_n3838_ = 1'b1;
3'b??1 : new_n3838_ = 1'b1;
default : new_n3838_ = 1'b0;
endcase
casez ({x[2], new_n290_, new_n294_})
3'b01? : new_n3839_ = 1'b1;
3'b??1 : new_n3839_ = 1'b1;
default : new_n3839_ = 1'b0;
endcase
casez ({new_n101_, new_n133_, new_n295_})
3'b11? : new_n3840_ = 1'b1;
3'b??1 : new_n3840_ = 1'b1;
default : new_n3840_ = 1'b0;
endcase
casez ({u[1], new_n243_, new_n295_})
3'b11? : new_n3841_ = 1'b1;
3'b??1 : new_n3841_ = 1'b1;
default : new_n3841_ = 1'b0;
endcase
casez ({new_n745_, new_n870_})
2'b00 : new_n3842_ = 1'b1;
default : new_n3842_ = 1'b0;
endcase
casez ({new_n107_, new_n206_, new_n295_})
3'b01? : new_n3843_ = 1'b1;
3'b??1 : new_n3843_ = 1'b1;
default : new_n3843_ = 1'b0;
endcase
casez ({u[2], new_n574_, new_n448_})
3'b10? : new_n3844_ = 1'b1;
3'b??1 : new_n3844_ = 1'b1;
default : new_n3844_ = 1'b0;
endcase
casez ({new_n448_, new_n871_})
2'b00 : new_n3845_ = 1'b1;
default : new_n3845_ = 1'b0;
endcase
casez ({new_n126_, new_n872_})
2'b00 : new_n3846_ = 1'b1;
default : new_n3846_ = 1'b0;
endcase
casez ({new_n321_, new_n439_, new_n577_})
3'b10? : new_n3847_ = 1'b1;
3'b??1 : new_n3847_ = 1'b1;
default : new_n3847_ = 1'b0;
endcase
casez ({new_n334_, new_n873_})
2'b00 : new_n3848_ = 1'b1;
default : new_n3848_ = 1'b0;
endcase
casez ({new_n378_, new_n1338_})
2'b00 : new_n3849_ = 1'b1;
default : new_n3849_ = 1'b0;
endcase
casez ({new_n162_, new_n285_, new_n1339_})
3'b11? : new_n3850_ = 1'b1;
3'b??1 : new_n3850_ = 1'b1;
default : new_n3850_ = 1'b0;
endcase
casez ({new_n290_, new_n578_})
2'b00 : new_n3851_ = 1'b1;
default : new_n3851_ = 1'b0;
endcase
casez ({u[1], new_n578_, new_n176_, new_n225_})
4'b11?? : new_n3852_ = 1'b1;
4'b??11 : new_n3852_ = 1'b1;
default : new_n3852_ = 1'b0;
endcase
casez ({new_n295_, new_n874_})
2'b00 : new_n3853_ = 1'b1;
default : new_n3853_ = 1'b0;
endcase
casez ({y[2], new_n336_, u[0], new_n579_})
4'b01?? : new_n3854_ = 1'b1;
4'b??01 : new_n3854_ = 1'b1;
default : new_n3854_ = 1'b0;
endcase
casez ({new_n1026_, new_n1340_})
2'b00 : new_n3855_ = 1'b1;
default : new_n3855_ = 1'b0;
endcase
casez ({new_n89_, new_n366_, new_n1340_})
3'b01? : new_n3856_ = 1'b1;
3'b??1 : new_n3856_ = 1'b1;
default : new_n3856_ = 1'b0;
endcase
casez ({new_n420_, new_n509_, new_n1341_})
3'b11? : new_n3857_ = 1'b1;
3'b??1 : new_n3857_ = 1'b1;
default : new_n3857_ = 1'b0;
endcase
casez ({new_n738_, new_n1341_})
2'b00 : new_n3858_ = 1'b1;
default : new_n3858_ = 1'b0;
endcase
casez ({new_n122_, new_n243_, new_n1341_})
3'b11? : new_n3859_ = 1'b1;
3'b??1 : new_n3859_ = 1'b1;
default : new_n3859_ = 1'b0;
endcase
casez ({x[1], new_n176_, new_n875_})
3'b11? : new_n3860_ = 1'b1;
3'b??1 : new_n3860_ = 1'b1;
default : new_n3860_ = 1'b0;
endcase
casez ({new_n93_, new_n176_, new_n875_})
3'b11? : new_n3861_ = 1'b1;
3'b??1 : new_n3861_ = 1'b1;
default : new_n3861_ = 1'b0;
endcase
casez ({new_n271_, new_n1343_})
2'b00 : new_n3862_ = 1'b1;
default : new_n3862_ = 1'b0;
endcase
casez ({new_n85_, new_n398_, new_n581_})
3'b11? : new_n3863_ = 1'b1;
3'b??1 : new_n3863_ = 1'b1;
default : new_n3863_ = 1'b0;
endcase
casez ({new_n677_, new_n1345_})
2'b00 : new_n3864_ = 1'b1;
default : new_n3864_ = 1'b0;
endcase
casez ({v[1], new_n324_, new_n1345_})
3'b01? : new_n3865_ = 1'b1;
3'b??1 : new_n3865_ = 1'b1;
default : new_n3865_ = 1'b0;
endcase
casez ({new_n4598_, new_n118_, new_n344_})
3'b1?? : new_n3866_ = 1'b1;
3'b?11 : new_n3866_ = 1'b1;
default : new_n3866_ = 1'b0;
endcase
casez ({new_n367_, new_n1347_})
2'b00 : new_n3867_ = 1'b1;
default : new_n3867_ = 1'b0;
endcase
casez ({new_n97_, new_n551_, new_n1347_})
3'b11? : new_n3868_ = 1'b1;
3'b??1 : new_n3868_ = 1'b1;
default : new_n3868_ = 1'b0;
endcase
casez ({new_n865_, new_n1349_})
2'b00 : new_n3869_ = 1'b1;
default : new_n3869_ = 1'b0;
endcase
casez ({new_n937_, new_n1349_})
2'b00 : new_n3870_ = 1'b1;
default : new_n3870_ = 1'b0;
endcase
casez ({new_n86_, new_n216_, new_n583_})
3'b11? : new_n3871_ = 1'b1;
3'b??1 : new_n3871_ = 1'b1;
default : new_n3871_ = 1'b0;
endcase
casez ({new_n310_, new_n583_})
2'b00 : new_n3872_ = 1'b1;
default : new_n3872_ = 1'b0;
endcase
casez ({new_n536_, new_n584_})
2'b00 : new_n3873_ = 1'b1;
default : new_n3873_ = 1'b0;
endcase
casez ({new_n525_, new_n584_})
2'b00 : new_n3874_ = 1'b1;
default : new_n3874_ = 1'b0;
endcase
casez ({new_n1114_, new_n1352_})
2'b00 : new_n3875_ = 1'b1;
default : new_n3875_ = 1'b0;
endcase
casez ({new_n4597_, new_n1353_})
2'b1? : new_n3876_ = 1'b1;
2'b?1 : new_n3876_ = 1'b1;
default : new_n3876_ = 1'b0;
endcase
casez ({new_n1346_, new_n1353_})
2'b00 : new_n3877_ = 1'b1;
default : new_n3877_ = 1'b0;
endcase
casez ({new_n244_, new_n619_, new_n1355_})
3'b11? : new_n3878_ = 1'b1;
3'b??1 : new_n3878_ = 1'b1;
default : new_n3878_ = 1'b0;
endcase
casez ({new_n129_, new_n508_, new_n1355_})
3'b11? : new_n3879_ = 1'b1;
3'b??1 : new_n3879_ = 1'b1;
default : new_n3879_ = 1'b0;
endcase
casez ({new_n738_, new_n1356_})
2'b00 : new_n3880_ = 1'b1;
default : new_n3880_ = 1'b0;
endcase
casez ({x[2], new_n1356_, new_n175_, new_n407_})
4'b11?? : new_n3881_ = 1'b1;
4'b??11 : new_n3881_ = 1'b1;
default : new_n3881_ = 1'b0;
endcase
casez ({new_n171_, new_n264_, new_n1356_})
3'b11? : new_n3882_ = 1'b1;
3'b??1 : new_n3882_ = 1'b1;
default : new_n3882_ = 1'b0;
endcase
casez ({new_n738_, new_n1357_})
2'b00 : new_n3883_ = 1'b1;
default : new_n3883_ = 1'b0;
endcase
casez ({new_n860_, new_n1358_})
2'b00 : new_n3884_ = 1'b1;
default : new_n3884_ = 1'b0;
endcase
casez ({new_n1015_, new_n1359_})
2'b00 : new_n3885_ = 1'b1;
default : new_n3885_ = 1'b0;
endcase
casez ({new_n160_, new_n241_, new_n1359_})
3'b11? : new_n3886_ = 1'b1;
3'b??1 : new_n3886_ = 1'b1;
default : new_n3886_ = 1'b0;
endcase
casez ({new_n118_, new_n933_, new_n1359_})
3'b10? : new_n3887_ = 1'b1;
3'b??1 : new_n3887_ = 1'b1;
default : new_n3887_ = 1'b0;
endcase
casez ({new_n295_, new_n1361_})
2'b00 : new_n3888_ = 1'b1;
default : new_n3888_ = 1'b0;
endcase
casez ({new_n857_, new_n1361_})
2'b00 : new_n3889_ = 1'b1;
default : new_n3889_ = 1'b0;
endcase
casez ({new_n80_, new_n89_, new_n1362_})
3'b11? : new_n3890_ = 1'b1;
3'b??1 : new_n3890_ = 1'b1;
default : new_n3890_ = 1'b0;
endcase
casez ({new_n1017_, new_n1365_})
2'b00 : new_n3891_ = 1'b1;
default : new_n3891_ = 1'b0;
endcase
casez ({y[2], new_n1129_, new_n1365_})
3'b01? : new_n3892_ = 1'b1;
3'b??1 : new_n3892_ = 1'b1;
default : new_n3892_ = 1'b0;
endcase
casez ({new_n638_, new_n1365_})
2'b00 : new_n3893_ = 1'b1;
default : new_n3893_ = 1'b0;
endcase
casez ({new_n1092_, new_n1366_})
2'b00 : new_n3894_ = 1'b1;
default : new_n3894_ = 1'b0;
endcase
casez ({new_n384_, new_n1368_})
2'b00 : new_n3895_ = 1'b1;
default : new_n3895_ = 1'b0;
endcase
casez ({new_n4646_, new_n1369_})
2'b1? : new_n3896_ = 1'b1;
2'b?1 : new_n3896_ = 1'b1;
default : new_n3896_ = 1'b0;
endcase
casez ({new_n639_, new_n1369_})
2'b00 : new_n3897_ = 1'b1;
default : new_n3897_ = 1'b0;
endcase
casez ({new_n1124_, new_n1369_})
2'b00 : new_n3898_ = 1'b1;
default : new_n3898_ = 1'b0;
endcase
casez ({new_n255_, new_n441_, new_n494_, new_n598_})
4'b11?? : new_n3899_ = 1'b1;
4'b??11 : new_n3899_ = 1'b1;
default : new_n3899_ = 1'b0;
endcase
casez ({new_n788_, new_n1369_})
2'b00 : new_n3900_ = 1'b1;
default : new_n3900_ = 1'b0;
endcase
casez ({new_n238_, new_n332_, new_n1371_})
3'b11? : new_n3901_ = 1'b1;
3'b??1 : new_n3901_ = 1'b1;
default : new_n3901_ = 1'b0;
endcase
casez ({new_n1030_, new_n1372_})
2'b00 : new_n3902_ = 1'b1;
default : new_n3902_ = 1'b0;
endcase
casez ({new_n127_, new_n430_, new_n1372_})
3'b11? : new_n3903_ = 1'b1;
3'b??1 : new_n3903_ = 1'b1;
default : new_n3903_ = 1'b0;
endcase
casez ({new_n121_, new_n131_, new_n600_})
3'b11? : new_n3904_ = 1'b1;
3'b??1 : new_n3904_ = 1'b1;
default : new_n3904_ = 1'b0;
endcase
casez ({new_n97_, new_n299_, new_n1373_})
3'b11? : new_n3905_ = 1'b1;
3'b??1 : new_n3905_ = 1'b1;
default : new_n3905_ = 1'b0;
endcase
casez ({new_n1105_, new_n1374_})
2'b00 : new_n3906_ = 1'b1;
default : new_n3906_ = 1'b0;
endcase
casez ({new_n151_, new_n218_, new_n1375_})
3'b11? : new_n3907_ = 1'b1;
3'b??1 : new_n3907_ = 1'b1;
default : new_n3907_ = 1'b0;
endcase
casez ({new_n396_, new_n478_, new_n601_})
3'b11? : new_n3908_ = 1'b1;
3'b??1 : new_n3908_ = 1'b1;
default : new_n3908_ = 1'b0;
endcase
casez ({new_n1154_, new_n1375_})
2'b00 : new_n3909_ = 1'b1;
default : new_n3909_ = 1'b0;
endcase
casez ({new_n103_, new_n495_, new_n601_})
3'b11? : new_n3910_ = 1'b1;
3'b??1 : new_n3910_ = 1'b1;
default : new_n3910_ = 1'b0;
endcase
casez ({new_n746_, new_n1376_})
2'b00 : new_n3911_ = 1'b1;
default : new_n3911_ = 1'b0;
endcase
casez ({u[1], new_n786_, new_n1377_})
3'b01? : new_n3912_ = 1'b1;
3'b??1 : new_n3912_ = 1'b1;
default : new_n3912_ = 1'b0;
endcase
casez ({new_n185_, new_n602_})
2'b00 : new_n3913_ = 1'b1;
default : new_n3913_ = 1'b0;
endcase
casez ({new_n79_, new_n308_, new_n602_})
3'b01? : new_n3914_ = 1'b1;
3'b??1 : new_n3914_ = 1'b1;
default : new_n3914_ = 1'b0;
endcase
casez ({v[2], new_n251_, new_n1377_})
3'b01? : new_n3915_ = 1'b1;
3'b??1 : new_n3915_ = 1'b1;
default : new_n3915_ = 1'b0;
endcase
casez ({x[1], new_n1378_, new_n1122_})
3'b11? : new_n3916_ = 1'b1;
3'b??1 : new_n3916_ = 1'b1;
default : new_n3916_ = 1'b0;
endcase
casez ({new_n89_, new_n181_, new_n602_})
3'b00? : new_n3917_ = 1'b1;
3'b??1 : new_n3917_ = 1'b1;
default : new_n3917_ = 1'b0;
endcase
casez ({new_n158_, new_n240_, new_n1380_})
3'b11? : new_n3918_ = 1'b1;
3'b??1 : new_n3918_ = 1'b1;
default : new_n3918_ = 1'b0;
endcase
casez ({new_n262_, new_n493_, new_n1381_})
3'b11? : new_n3919_ = 1'b1;
3'b??1 : new_n3919_ = 1'b1;
default : new_n3919_ = 1'b0;
endcase
casez ({new_n620_, new_n1383_})
2'b00 : new_n3920_ = 1'b1;
default : new_n3920_ = 1'b0;
endcase
casez ({x[1], new_n484_, new_n343_, new_n606_})
4'b11?? : new_n3921_ = 1'b1;
4'b??11 : new_n3921_ = 1'b1;
default : new_n3921_ = 1'b0;
endcase
casez ({new_n779_, new_n1383_})
2'b00 : new_n3922_ = 1'b1;
default : new_n3922_ = 1'b0;
endcase
casez ({new_n84_, new_n554_, new_n1384_})
3'b11? : new_n3923_ = 1'b1;
3'b??1 : new_n3923_ = 1'b1;
default : new_n3923_ = 1'b0;
endcase
casez ({new_n89_, new_n335_, new_n1384_})
3'b01? : new_n3924_ = 1'b1;
3'b??1 : new_n3924_ = 1'b1;
default : new_n3924_ = 1'b0;
endcase
casez ({new_n171_, new_n1047_, new_n225_, new_n1385_})
4'b11?? : new_n3925_ = 1'b1;
4'b??11 : new_n3925_ = 1'b1;
default : new_n3925_ = 1'b0;
endcase
casez ({new_n749_, new_n1385_})
2'b00 : new_n3926_ = 1'b1;
default : new_n3926_ = 1'b0;
endcase
casez ({new_n634_, new_n1386_})
2'b00 : new_n3927_ = 1'b1;
default : new_n3927_ = 1'b0;
endcase
casez ({new_n493_, new_n606_, new_n605_, new_n2498_})
4'b11?? : new_n3928_ = 1'b1;
4'b??11 : new_n3928_ = 1'b1;
default : new_n3928_ = 1'b0;
endcase
casez ({new_n669_, new_n1388_})
2'b00 : new_n3929_ = 1'b1;
default : new_n3929_ = 1'b0;
endcase
casez ({new_n161_, new_n417_, new_n1389_})
3'b11? : new_n3930_ = 1'b1;
3'b??1 : new_n3930_ = 1'b1;
default : new_n3930_ = 1'b0;
endcase
casez ({new_n1172_, new_n1389_})
2'b00 : new_n3931_ = 1'b1;
default : new_n3931_ = 1'b0;
endcase
casez ({x[2], new_n169_, new_n1389_})
3'b11? : new_n3932_ = 1'b1;
3'b??1 : new_n3932_ = 1'b1;
default : new_n3932_ = 1'b0;
endcase
casez ({new_n225_, new_n579_, new_n320_, new_n1390_})
4'b11?? : new_n3933_ = 1'b1;
4'b??01 : new_n3933_ = 1'b1;
default : new_n3933_ = 1'b0;
endcase
casez ({new_n1100_, new_n2511_})
2'b10 : new_n3934_ = 1'b1;
default : new_n3934_ = 1'b0;
endcase
casez ({new_n1016_, new_n2516_})
2'b00 : new_n3935_ = 1'b1;
default : new_n3935_ = 1'b0;
endcase
casez ({new_n441_, new_n1392_})
2'b00 : new_n3936_ = 1'b1;
default : new_n3936_ = 1'b0;
endcase
casez ({new_n239_, new_n496_, new_n350_, new_n2518_})
4'b11?? : new_n3937_ = 1'b1;
4'b??11 : new_n3937_ = 1'b1;
default : new_n3937_ = 1'b0;
endcase
casez ({new_n207_, new_n2523_, new_n1934_})
3'b10? : new_n3938_ = 1'b1;
3'b??1 : new_n3938_ = 1'b1;
default : new_n3938_ = 1'b0;
endcase
casez ({new_n224_, new_n2525_, new_n1869_})
3'b10? : new_n3939_ = 1'b1;
3'b??1 : new_n3939_ = 1'b1;
default : new_n3939_ = 1'b0;
endcase
casez ({new_n198_, new_n2527_, new_n1887_})
3'b10? : new_n3940_ = 1'b1;
3'b??1 : new_n3940_ = 1'b1;
default : new_n3940_ = 1'b0;
endcase
casez ({new_n308_, new_n654_, new_n456_, new_n2531_})
4'b11?? : new_n3941_ = 1'b1;
4'b??10 : new_n3941_ = 1'b1;
default : new_n3941_ = 1'b0;
endcase
casez ({new_n131_, new_n2532_, new_n1836_})
3'b10? : new_n3942_ = 1'b1;
3'b??1 : new_n3942_ = 1'b1;
default : new_n3942_ = 1'b0;
endcase
casez ({new_n151_, new_n2533_, new_n1609_})
3'b10? : new_n3943_ = 1'b1;
3'b??1 : new_n3943_ = 1'b1;
default : new_n3943_ = 1'b0;
endcase
casez ({new_n249_, new_n1035_, new_n381_, new_n2535_})
4'b11?? : new_n3944_ = 1'b1;
4'b??10 : new_n3944_ = 1'b1;
default : new_n3944_ = 1'b0;
endcase
casez ({new_n92_, new_n2536_, new_n857_})
3'b10? : new_n3945_ = 1'b1;
3'b??1 : new_n3945_ = 1'b1;
default : new_n3945_ = 1'b0;
endcase
casez ({y[2], new_n2537_, new_n962_})
3'b00? : new_n3946_ = 1'b1;
3'b??1 : new_n3946_ = 1'b1;
default : new_n3946_ = 1'b0;
endcase
casez ({new_n142_, new_n2545_, new_n169_, new_n2544_})
4'b10?? : new_n3947_ = 1'b1;
4'b??10 : new_n3947_ = 1'b1;
default : new_n3947_ = 1'b0;
endcase
casez ({new_n162_, new_n439_, new_n321_, new_n2548_})
4'b10?? : new_n3948_ = 1'b1;
4'b??10 : new_n3948_ = 1'b1;
default : new_n3948_ = 1'b0;
endcase
casez ({u[0], new_n2550_, new_n239_})
3'b00? : new_n3949_ = 1'b1;
3'b??1 : new_n3949_ = 1'b1;
default : new_n3949_ = 1'b0;
endcase
casez ({y[2], new_n2553_, new_n539_})
3'b11? : new_n3950_ = 1'b1;
3'b??1 : new_n3950_ = 1'b1;
default : new_n3950_ = 1'b0;
endcase
casez ({new_n148_, new_n2553_, new_n157_, new_n162_})
4'b11?? : new_n3951_ = 1'b1;
4'b??11 : new_n3951_ = 1'b1;
default : new_n3951_ = 1'b0;
endcase
casez ({new_n384_, new_n2554_})
2'b00 : new_n3952_ = 1'b1;
default : new_n3952_ = 1'b0;
endcase
casez ({new_n4585_, new_n2554_})
2'b1? : new_n3953_ = 1'b1;
2'b?1 : new_n3953_ = 1'b1;
default : new_n3953_ = 1'b0;
endcase
casez ({new_n4599_, new_n280_})
2'b1? : new_n3954_ = 1'b1;
2'b?1 : new_n3954_ = 1'b1;
default : new_n3954_ = 1'b0;
endcase
casez ({new_n303_, new_n1394_})
2'b00 : new_n3955_ = 1'b1;
default : new_n3955_ = 1'b0;
endcase
casez ({new_n129_, new_n444_, new_n2558_})
3'b11? : new_n3956_ = 1'b1;
3'b??1 : new_n3956_ = 1'b1;
default : new_n3956_ = 1'b0;
endcase
casez ({new_n858_, new_n2559_})
2'b00 : new_n3957_ = 1'b1;
default : new_n3957_ = 1'b0;
endcase
casez ({new_n89_, new_n1570_, new_n2559_})
3'b11? : new_n3958_ = 1'b1;
3'b??1 : new_n3958_ = 1'b1;
default : new_n3958_ = 1'b0;
endcase
casez ({new_n1831_, new_n2560_})
2'b00 : new_n3959_ = 1'b1;
default : new_n3959_ = 1'b0;
endcase
casez ({new_n1042_, new_n1395_})
2'b00 : new_n3960_ = 1'b1;
default : new_n3960_ = 1'b0;
endcase
casez ({new_n1162_, new_n1396_})
2'b00 : new_n3961_ = 1'b1;
default : new_n3961_ = 1'b0;
endcase
casez ({new_n1560_, new_n2562_})
2'b00 : new_n3962_ = 1'b1;
default : new_n3962_ = 1'b0;
endcase
casez ({new_n278_, new_n369_, new_n1396_})
3'b11? : new_n3963_ = 1'b1;
3'b??1 : new_n3963_ = 1'b1;
default : new_n3963_ = 1'b0;
endcase
casez ({new_n1364_, new_n2562_})
2'b00 : new_n3964_ = 1'b1;
default : new_n3964_ = 1'b0;
endcase
casez ({new_n4630_, new_n2562_})
2'b1? : new_n3965_ = 1'b1;
2'b?1 : new_n3965_ = 1'b1;
default : new_n3965_ = 1'b0;
endcase
casez ({new_n424_, new_n1396_})
2'b00 : new_n3966_ = 1'b1;
default : new_n3966_ = 1'b0;
endcase
casez ({new_n675_, new_n1396_})
2'b00 : new_n3967_ = 1'b1;
default : new_n3967_ = 1'b0;
endcase
casez ({new_n1393_, new_n1397_})
2'b00 : new_n3968_ = 1'b1;
default : new_n3968_ = 1'b0;
endcase
casez ({new_n873_, new_n1397_})
2'b00 : new_n3969_ = 1'b1;
default : new_n3969_ = 1'b0;
endcase
casez ({u[2], new_n259_, new_n2568_})
3'b11? : new_n3970_ = 1'b1;
3'b??1 : new_n3970_ = 1'b1;
default : new_n3970_ = 1'b0;
endcase
casez ({new_n1582_, new_n2568_})
2'b00 : new_n3971_ = 1'b1;
default : new_n3971_ = 1'b0;
endcase
casez ({new_n1008_, new_n2569_})
2'b00 : new_n3972_ = 1'b1;
default : new_n3972_ = 1'b0;
endcase
casez ({new_n259_, new_n1399_})
2'b00 : new_n3973_ = 1'b1;
default : new_n3973_ = 1'b0;
endcase
casez ({new_n1391_, new_n2571_})
2'b00 : new_n3974_ = 1'b1;
default : new_n3974_ = 1'b0;
endcase
casez ({new_n636_, new_n1400_})
2'b00 : new_n3975_ = 1'b1;
default : new_n3975_ = 1'b0;
endcase
casez ({new_n407_, new_n2573_})
2'b00 : new_n3976_ = 1'b1;
default : new_n3976_ = 1'b0;
endcase
casez ({new_n1608_, new_n2573_})
2'b00 : new_n3977_ = 1'b1;
default : new_n3977_ = 1'b0;
endcase
casez ({new_n83_, new_n1401_, new_n84_, new_n448_})
4'b11?? : new_n3978_ = 1'b1;
4'b??11 : new_n3978_ = 1'b1;
default : new_n3978_ = 1'b0;
endcase
casez ({new_n1039_, new_n1401_})
2'b00 : new_n3979_ = 1'b1;
default : new_n3979_ = 1'b0;
endcase
casez ({new_n79_, new_n1002_, new_n2575_})
3'b11? : new_n3980_ = 1'b1;
3'b??1 : new_n3980_ = 1'b1;
default : new_n3980_ = 1'b0;
endcase
casez ({x[1], new_n133_, new_n1402_})
3'b01? : new_n3981_ = 1'b1;
3'b??1 : new_n3981_ = 1'b1;
default : new_n3981_ = 1'b0;
endcase
casez ({new_n1596_, new_n2576_})
2'b00 : new_n3982_ = 1'b1;
default : new_n3982_ = 1'b0;
endcase
casez ({new_n1839_, new_n2576_})
2'b00 : new_n3983_ = 1'b1;
default : new_n3983_ = 1'b0;
endcase
casez ({new_n455_, new_n1402_})
2'b00 : new_n3984_ = 1'b1;
default : new_n3984_ = 1'b0;
endcase
casez ({new_n1373_, new_n1403_})
2'b00 : new_n3985_ = 1'b1;
default : new_n3985_ = 1'b0;
endcase
casez ({new_n404_, new_n2579_})
2'b00 : new_n3986_ = 1'b1;
default : new_n3986_ = 1'b0;
endcase
casez ({new_n1857_, new_n2580_})
2'b00 : new_n3987_ = 1'b1;
default : new_n3987_ = 1'b0;
endcase
casez ({new_n870_, new_n2580_})
2'b00 : new_n3988_ = 1'b1;
default : new_n3988_ = 1'b0;
endcase
casez ({new_n775_, new_n2581_})
2'b00 : new_n3989_ = 1'b1;
default : new_n3989_ = 1'b0;
endcase
casez ({new_n1939_, new_n2584_})
2'b00 : new_n3990_ = 1'b1;
default : new_n3990_ = 1'b0;
endcase
casez ({new_n777_, new_n2585_})
2'b00 : new_n3991_ = 1'b1;
default : new_n3991_ = 1'b0;
endcase
casez ({new_n2556_, new_n2586_})
2'b00 : new_n3992_ = 1'b1;
default : new_n3992_ = 1'b0;
endcase
casez ({new_n631_, new_n2588_})
2'b00 : new_n3993_ = 1'b1;
default : new_n3993_ = 1'b0;
endcase
casez ({new_n2560_, new_n2589_})
2'b00 : new_n3994_ = 1'b1;
default : new_n3994_ = 1'b0;
endcase
casez ({new_n1371_, new_n2590_})
2'b00 : new_n3995_ = 1'b1;
default : new_n3995_ = 1'b0;
endcase
casez ({x[1], new_n557_, new_n617_})
3'b01? : new_n3996_ = 1'b1;
3'b??1 : new_n3996_ = 1'b1;
default : new_n3996_ = 1'b0;
endcase
casez ({new_n347_, new_n2592_})
2'b00 : new_n3997_ = 1'b1;
default : new_n3997_ = 1'b0;
endcase
casez ({new_n635_, new_n2592_})
2'b00 : new_n3998_ = 1'b1;
default : new_n3998_ = 1'b0;
endcase
casez ({new_n142_, new_n178_, new_n2595_})
3'b11? : new_n3999_ = 1'b1;
3'b??1 : new_n3999_ = 1'b1;
default : new_n3999_ = 1'b0;
endcase
casez ({new_n1905_, new_n2596_})
2'b00 : new_n4000_ = 1'b1;
default : new_n4000_ = 1'b0;
endcase
casez ({new_n1044_, new_n2597_})
2'b00 : new_n4001_ = 1'b1;
default : new_n4001_ = 1'b0;
endcase
casez ({new_n1874_, new_n2597_})
2'b00 : new_n4002_ = 1'b1;
default : new_n4002_ = 1'b0;
endcase
casez ({new_n857_, new_n2598_})
2'b00 : new_n4003_ = 1'b1;
default : new_n4003_ = 1'b0;
endcase
casez ({new_n4621_, new_n2598_})
2'b1? : new_n4004_ = 1'b1;
2'b?1 : new_n4004_ = 1'b1;
default : new_n4004_ = 1'b0;
endcase
casez ({new_n1856_, new_n2600_})
2'b00 : new_n4005_ = 1'b1;
default : new_n4005_ = 1'b0;
endcase
casez ({new_n1612_, new_n2600_})
2'b00 : new_n4006_ = 1'b1;
default : new_n4006_ = 1'b0;
endcase
casez ({new_n581_, new_n2600_})
2'b00 : new_n4007_ = 1'b1;
default : new_n4007_ = 1'b0;
endcase
casez ({new_n83_, new_n347_, new_n2601_})
3'b11? : new_n4008_ = 1'b1;
3'b??1 : new_n4008_ = 1'b1;
default : new_n4008_ = 1'b0;
endcase
casez ({new_n1618_, new_n2601_})
2'b00 : new_n4009_ = 1'b1;
default : new_n4009_ = 1'b0;
endcase
casez ({new_n369_, new_n2546_, new_n2602_})
3'b10? : new_n4010_ = 1'b1;
3'b??1 : new_n4010_ = 1'b1;
default : new_n4010_ = 1'b0;
endcase
casez ({new_n1122_, new_n2603_})
2'b00 : new_n4011_ = 1'b1;
default : new_n4011_ = 1'b0;
endcase
casez ({new_n267_, new_n924_})
2'b00 : new_n4012_ = 1'b1;
default : new_n4012_ = 1'b0;
endcase
casez ({new_n83_, new_n558_, new_n198_, new_n925_})
4'b01?? : new_n4013_ = 1'b1;
4'b??10 : new_n4013_ = 1'b1;
default : new_n4013_ = 1'b0;
endcase
casez ({new_n95_, new_n925_, new_n632_})
3'b10? : new_n4014_ = 1'b1;
3'b??1 : new_n4014_ = 1'b1;
default : new_n4014_ = 1'b0;
endcase
casez ({new_n202_, new_n618_})
2'b00 : new_n4015_ = 1'b1;
default : new_n4015_ = 1'b0;
endcase
casez ({new_n317_, new_n394_, new_n2604_})
3'b10? : new_n4016_ = 1'b1;
3'b??1 : new_n4016_ = 1'b1;
default : new_n4016_ = 1'b0;
endcase
casez ({new_n1927_, new_n2605_})
2'b00 : new_n4017_ = 1'b1;
default : new_n4017_ = 1'b0;
endcase
casez ({new_n1611_, new_n2606_})
2'b00 : new_n4018_ = 1'b1;
default : new_n4018_ = 1'b0;
endcase
casez ({new_n1918_, new_n2607_})
2'b00 : new_n4019_ = 1'b1;
default : new_n4019_ = 1'b0;
endcase
casez ({new_n140_, new_n186_})
2'b00 : new_n4020_ = 1'b1;
default : new_n4020_ = 1'b0;
endcase
casez ({new_n91_, new_n398_, new_n598_, new_n619_})
4'b11?? : new_n4021_ = 1'b1;
4'b??11 : new_n4021_ = 1'b1;
default : new_n4021_ = 1'b0;
endcase
casez ({new_n2606_, new_n2609_})
2'b00 : new_n4022_ = 1'b1;
default : new_n4022_ = 1'b0;
endcase
casez ({new_n945_, new_n2609_})
2'b00 : new_n4023_ = 1'b1;
default : new_n4023_ = 1'b0;
endcase
casez ({new_n231_, new_n250_, new_n2610_})
3'b11? : new_n4024_ = 1'b1;
3'b??1 : new_n4024_ = 1'b1;
default : new_n4024_ = 1'b0;
endcase
casez ({new_n535_, new_n2610_})
2'b00 : new_n4025_ = 1'b1;
default : new_n4025_ = 1'b0;
endcase
casez ({new_n169_, new_n933_, new_n384_})
3'b10? : new_n4026_ = 1'b1;
3'b??1 : new_n4026_ = 1'b1;
default : new_n4026_ = 1'b0;
endcase
casez ({new_n1595_, new_n2613_})
2'b00 : new_n4027_ = 1'b1;
default : new_n4027_ = 1'b0;
endcase
casez ({new_n208_, new_n332_, new_n2613_})
3'b11? : new_n4028_ = 1'b1;
3'b??1 : new_n4028_ = 1'b1;
default : new_n4028_ = 1'b0;
endcase
casez ({new_n1838_, new_n2614_})
2'b00 : new_n4029_ = 1'b1;
default : new_n4029_ = 1'b0;
endcase
casez ({new_n1588_, new_n2614_})
2'b00 : new_n4030_ = 1'b1;
default : new_n4030_ = 1'b0;
endcase
casez ({new_n1920_, new_n2615_})
2'b00 : new_n4031_ = 1'b1;
default : new_n4031_ = 1'b0;
endcase
casez ({new_n2585_, new_n2616_})
2'b00 : new_n4032_ = 1'b1;
default : new_n4032_ = 1'b0;
endcase
casez ({new_n150_, new_n1544_, new_n2616_})
3'b11? : new_n4033_ = 1'b1;
3'b??1 : new_n4033_ = 1'b1;
default : new_n4033_ = 1'b0;
endcase
casez ({new_n1388_, new_n2617_})
2'b00 : new_n4034_ = 1'b1;
default : new_n4034_ = 1'b0;
endcase
casez ({new_n1645_, new_n2617_})
2'b00 : new_n4035_ = 1'b1;
default : new_n4035_ = 1'b0;
endcase
casez ({new_n740_, new_n2618_})
2'b00 : new_n4036_ = 1'b1;
default : new_n4036_ = 1'b0;
endcase
casez ({new_n151_, new_n250_, new_n2618_})
3'b11? : new_n4037_ = 1'b1;
3'b??1 : new_n4037_ = 1'b1;
default : new_n4037_ = 1'b0;
endcase
casez ({new_n268_, new_n2620_})
2'b00 : new_n4038_ = 1'b1;
default : new_n4038_ = 1'b0;
endcase
casez ({new_n334_, new_n2620_})
2'b00 : new_n4039_ = 1'b1;
default : new_n4039_ = 1'b0;
endcase
casez ({new_n1917_, new_n2621_})
2'b00 : new_n4040_ = 1'b1;
default : new_n4040_ = 1'b0;
endcase
casez ({new_n1946_, new_n2621_})
2'b00 : new_n4041_ = 1'b1;
default : new_n4041_ = 1'b0;
endcase
casez ({new_n251_, new_n2621_})
2'b00 : new_n4042_ = 1'b1;
default : new_n4042_ = 1'b0;
endcase
casez ({new_n1586_, new_n2622_})
2'b00 : new_n4043_ = 1'b1;
default : new_n4043_ = 1'b0;
endcase
casez ({new_n101_, new_n340_, new_n2623_})
3'b01? : new_n4044_ = 1'b1;
3'b??1 : new_n4044_ = 1'b1;
default : new_n4044_ = 1'b0;
endcase
casez ({new_n290_, new_n2624_})
2'b00 : new_n4045_ = 1'b1;
default : new_n4045_ = 1'b0;
endcase
casez ({x[2], new_n271_, new_n2624_})
3'b11? : new_n4046_ = 1'b1;
3'b??1 : new_n4046_ = 1'b1;
default : new_n4046_ = 1'b0;
endcase
casez ({y[1], new_n483_, new_n2624_})
3'b01? : new_n4047_ = 1'b1;
3'b??1 : new_n4047_ = 1'b1;
default : new_n4047_ = 1'b0;
endcase
casez ({new_n190_, new_n2625_})
2'b00 : new_n4048_ = 1'b1;
default : new_n4048_ = 1'b0;
endcase
casez ({new_n1565_, new_n2626_})
2'b00 : new_n4049_ = 1'b1;
default : new_n4049_ = 1'b0;
endcase
casez ({new_n419_, new_n2627_})
2'b00 : new_n4050_ = 1'b1;
default : new_n4050_ = 1'b0;
endcase
casez ({new_n161_, new_n509_, new_n2627_})
3'b11? : new_n4051_ = 1'b1;
3'b??1 : new_n4051_ = 1'b1;
default : new_n4051_ = 1'b0;
endcase
casez ({new_n857_, new_n939_})
2'b00 : new_n4052_ = 1'b1;
default : new_n4052_ = 1'b0;
endcase
casez ({new_n184_, new_n264_, new_n2628_})
3'b11? : new_n4053_ = 1'b1;
3'b??1 : new_n4053_ = 1'b1;
default : new_n4053_ = 1'b0;
endcase
casez ({new_n540_, new_n939_})
2'b00 : new_n4054_ = 1'b1;
default : new_n4054_ = 1'b0;
endcase
casez ({new_n1560_, new_n2629_})
2'b00 : new_n4055_ = 1'b1;
default : new_n4055_ = 1'b0;
endcase
casez ({new_n2602_, new_n2629_})
2'b00 : new_n4056_ = 1'b1;
default : new_n4056_ = 1'b0;
endcase
casez ({new_n955_, new_n2630_})
2'b00 : new_n4057_ = 1'b1;
default : new_n4057_ = 1'b0;
endcase
casez ({new_n743_, new_n2630_})
2'b00 : new_n4058_ = 1'b1;
default : new_n4058_ = 1'b0;
endcase
casez ({new_n737_, new_n2631_})
2'b00 : new_n4059_ = 1'b1;
default : new_n4059_ = 1'b0;
endcase
casez ({new_n1608_, new_n2631_})
2'b00 : new_n4060_ = 1'b1;
default : new_n4060_ = 1'b0;
endcase
casez ({new_n552_, new_n940_})
2'b00 : new_n4061_ = 1'b1;
default : new_n4061_ = 1'b0;
endcase
casez ({new_n745_, new_n2633_})
2'b00 : new_n4062_ = 1'b1;
default : new_n4062_ = 1'b0;
endcase
casez ({x[0], new_n109_, new_n206_, new_n2636_})
4'b001? : new_n4063_ = 1'b1;
4'b???1 : new_n4063_ = 1'b1;
default : new_n4063_ = 1'b0;
endcase
casez ({new_n1572_, new_n2636_})
2'b00 : new_n4064_ = 1'b1;
default : new_n4064_ = 1'b0;
endcase
casez ({new_n1576_, new_n2637_})
2'b00 : new_n4065_ = 1'b1;
default : new_n4065_ = 1'b0;
endcase
casez ({new_n4602_, new_n581_})
2'b1? : new_n4066_ = 1'b1;
2'b?1 : new_n4066_ = 1'b1;
default : new_n4066_ = 1'b0;
endcase
casez ({new_n4602_, new_n79_, new_n1178_})
3'b1?? : new_n4067_ = 1'b1;
3'b?01 : new_n4067_ = 1'b1;
default : new_n4067_ = 1'b0;
endcase
casez ({new_n2626_, new_n2640_})
2'b00 : new_n4068_ = 1'b1;
default : new_n4068_ = 1'b0;
endcase
casez ({new_n1118_, new_n2640_})
2'b00 : new_n4069_ = 1'b1;
default : new_n4069_ = 1'b0;
endcase
casez ({new_n1138_, new_n2641_})
2'b00 : new_n4070_ = 1'b1;
default : new_n4070_ = 1'b0;
endcase
casez ({new_n4614_, new_n2642_})
2'b1? : new_n4071_ = 1'b1;
2'b?1 : new_n4071_ = 1'b1;
default : new_n4071_ = 1'b0;
endcase
casez ({new_n543_, new_n941_})
2'b00 : new_n4072_ = 1'b1;
default : new_n4072_ = 1'b0;
endcase
casez ({new_n1894_, new_n2644_})
2'b00 : new_n4073_ = 1'b1;
default : new_n4073_ = 1'b0;
endcase
casez ({new_n729_, new_n941_})
2'b00 : new_n4074_ = 1'b1;
default : new_n4074_ = 1'b0;
endcase
casez ({v[2], new_n287_, new_n766_, new_n2645_})
4'b111? : new_n4075_ = 1'b1;
4'b???1 : new_n4075_ = 1'b1;
default : new_n4075_ = 1'b0;
endcase
casez ({u[0], new_n382_, new_n2645_})
3'b01? : new_n4076_ = 1'b1;
3'b??1 : new_n4076_ = 1'b1;
default : new_n4076_ = 1'b0;
endcase
casez ({new_n1856_, new_n2647_})
2'b00 : new_n4077_ = 1'b1;
default : new_n4077_ = 1'b0;
endcase
casez ({new_n1152_, new_n2648_})
2'b00 : new_n4078_ = 1'b1;
default : new_n4078_ = 1'b0;
endcase
casez ({new_n862_, new_n2650_})
2'b00 : new_n4079_ = 1'b1;
default : new_n4079_ = 1'b0;
endcase
casez ({new_n1916_, new_n2658_})
2'b00 : new_n4080_ = 1'b1;
default : new_n4080_ = 1'b0;
endcase
casez ({new_n1017_, new_n2658_})
2'b00 : new_n4081_ = 1'b1;
default : new_n4081_ = 1'b0;
endcase
casez ({new_n103_, new_n411_, new_n2658_})
3'b11? : new_n4082_ = 1'b1;
3'b??1 : new_n4082_ = 1'b1;
default : new_n4082_ = 1'b0;
endcase
casez ({new_n1149_, new_n2659_})
2'b00 : new_n4083_ = 1'b1;
default : new_n4083_ = 1'b0;
endcase
casez ({new_n1854_, new_n2660_})
2'b00 : new_n4084_ = 1'b1;
default : new_n4084_ = 1'b0;
endcase
casez ({new_n954_, new_n2660_})
2'b00 : new_n4085_ = 1'b1;
default : new_n4085_ = 1'b0;
endcase
casez ({new_n4601_, new_n2662_})
2'b1? : new_n4086_ = 1'b1;
2'b?1 : new_n4086_ = 1'b1;
default : new_n4086_ = 1'b0;
endcase
casez ({new_n4598_, new_n944_})
2'b1? : new_n4087_ = 1'b1;
2'b?1 : new_n4087_ = 1'b1;
default : new_n4087_ = 1'b0;
endcase
casez ({new_n419_, new_n2662_})
2'b00 : new_n4088_ = 1'b1;
default : new_n4088_ = 1'b0;
endcase
casez ({new_n1602_, new_n2664_})
2'b00 : new_n4089_ = 1'b1;
default : new_n4089_ = 1'b0;
endcase
casez ({new_n1115_, new_n2665_})
2'b00 : new_n4090_ = 1'b1;
default : new_n4090_ = 1'b0;
endcase
casez ({new_n471_, new_n2665_})
2'b00 : new_n4091_ = 1'b1;
default : new_n4091_ = 1'b0;
endcase
casez ({new_n121_, new_n196_, new_n2668_})
3'b11? : new_n4092_ = 1'b1;
3'b??1 : new_n4092_ = 1'b1;
default : new_n4092_ = 1'b0;
endcase
casez ({new_n103_, new_n616_, new_n2669_})
3'b11? : new_n4093_ = 1'b1;
3'b??1 : new_n4093_ = 1'b1;
default : new_n4093_ = 1'b0;
endcase
casez ({new_n718_, new_n2669_})
2'b00 : new_n4094_ = 1'b1;
default : new_n4094_ = 1'b0;
endcase
casez ({new_n2578_, new_n2672_})
2'b00 : new_n4095_ = 1'b1;
default : new_n4095_ = 1'b0;
endcase
casez ({new_n210_, new_n341_, new_n222_, new_n628_})
4'b11?? : new_n4096_ = 1'b1;
4'b??10 : new_n4096_ = 1'b1;
default : new_n4096_ = 1'b0;
endcase
casez ({new_n451_, new_n946_})
2'b00 : new_n4097_ = 1'b1;
default : new_n4097_ = 1'b0;
endcase
casez ({new_n1030_, new_n2674_})
2'b00 : new_n4098_ = 1'b1;
default : new_n4098_ = 1'b0;
endcase
casez ({new_n944_, new_n946_})
2'b00 : new_n4099_ = 1'b1;
default : new_n4099_ = 1'b0;
endcase
casez ({new_n1573_, new_n2675_})
2'b00 : new_n4100_ = 1'b1;
default : new_n4100_ = 1'b0;
endcase
casez ({new_n456_, new_n2678_})
2'b00 : new_n4101_ = 1'b1;
default : new_n4101_ = 1'b0;
endcase
casez ({new_n1019_, new_n2678_})
2'b00 : new_n4102_ = 1'b1;
default : new_n4102_ = 1'b0;
endcase
casez ({new_n207_, new_n439_, new_n2679_})
3'b10? : new_n4103_ = 1'b1;
3'b??1 : new_n4103_ = 1'b1;
default : new_n4103_ = 1'b0;
endcase
casez ({new_n775_, new_n2679_})
2'b00 : new_n4104_ = 1'b1;
default : new_n4104_ = 1'b0;
endcase
casez ({new_n274_, new_n998_, new_n2680_})
3'b10? : new_n4105_ = 1'b1;
3'b??1 : new_n4105_ = 1'b1;
default : new_n4105_ = 1'b0;
endcase
casez ({new_n2650_, new_n2681_})
2'b00 : new_n4106_ = 1'b1;
default : new_n4106_ = 1'b0;
endcase
casez ({new_n718_, new_n2682_})
2'b00 : new_n4107_ = 1'b1;
default : new_n4107_ = 1'b0;
endcase
casez ({new_n785_, new_n2682_})
2'b00 : new_n4108_ = 1'b1;
default : new_n4108_ = 1'b0;
endcase
casez ({y[2], new_n530_, new_n2685_})
3'b11? : new_n4109_ = 1'b1;
3'b??1 : new_n4109_ = 1'b1;
default : new_n4109_ = 1'b0;
endcase
casez ({new_n1114_, new_n2686_})
2'b00 : new_n4110_ = 1'b1;
default : new_n4110_ = 1'b0;
endcase
casez ({new_n4659_, new_n2688_})
2'b1? : new_n4111_ = 1'b1;
2'b?1 : new_n4111_ = 1'b1;
default : new_n4111_ = 1'b0;
endcase
casez ({new_n1109_, new_n2691_})
2'b00 : new_n4112_ = 1'b1;
default : new_n4112_ = 1'b0;
endcase
casez ({new_n944_, new_n2692_})
2'b00 : new_n4113_ = 1'b1;
default : new_n4113_ = 1'b0;
endcase
casez ({new_n4593_, new_n631_})
2'b1? : new_n4114_ = 1'b1;
2'b?1 : new_n4114_ = 1'b1;
default : new_n4114_ = 1'b0;
endcase
casez ({new_n1847_, new_n2693_})
2'b00 : new_n4115_ = 1'b1;
default : new_n4115_ = 1'b0;
endcase
casez ({new_n1895_, new_n2693_})
2'b00 : new_n4116_ = 1'b1;
default : new_n4116_ = 1'b0;
endcase
casez ({new_n797_, new_n2695_})
2'b00 : new_n4117_ = 1'b1;
default : new_n4117_ = 1'b0;
endcase
casez ({new_n940_, new_n2695_})
2'b00 : new_n4118_ = 1'b1;
default : new_n4118_ = 1'b0;
endcase
casez ({new_n4603_, new_n578_})
2'b1? : new_n4119_ = 1'b1;
2'b?1 : new_n4119_ = 1'b1;
default : new_n4119_ = 1'b0;
endcase
casez ({y[2], new_n2534_, new_n2697_})
3'b00? : new_n4120_ = 1'b1;
3'b??1 : new_n4120_ = 1'b1;
default : new_n4120_ = 1'b0;
endcase
casez ({new_n4603_, new_n601_})
2'b1? : new_n4121_ = 1'b1;
2'b?1 : new_n4121_ = 1'b1;
default : new_n4121_ = 1'b0;
endcase
casez ({new_n367_, new_n2698_})
2'b00 : new_n4122_ = 1'b1;
default : new_n4122_ = 1'b0;
endcase
casez ({new_n1353_, new_n2699_})
2'b00 : new_n4123_ = 1'b1;
default : new_n4123_ = 1'b0;
endcase
casez ({new_n1010_, new_n2699_})
2'b00 : new_n4124_ = 1'b1;
default : new_n4124_ = 1'b0;
endcase
casez ({x[0], new_n335_, new_n2699_})
3'b01? : new_n4125_ = 1'b1;
3'b??1 : new_n4125_ = 1'b1;
default : new_n4125_ = 1'b0;
endcase
casez ({new_n1634_, new_n2700_})
2'b00 : new_n4126_ = 1'b1;
default : new_n4126_ = 1'b0;
endcase
casez ({new_n738_, new_n2701_})
2'b00 : new_n4127_ = 1'b1;
default : new_n4127_ = 1'b0;
endcase
casez ({new_n1572_, new_n2702_})
2'b00 : new_n4128_ = 1'b1;
default : new_n4128_ = 1'b0;
endcase
casez ({new_n284_, new_n961_, new_n2703_})
3'b11? : new_n4129_ = 1'b1;
3'b??1 : new_n4129_ = 1'b1;
default : new_n4129_ = 1'b0;
endcase
casez ({new_n631_, new_n949_})
2'b00 : new_n4130_ = 1'b1;
default : new_n4130_ = 1'b0;
endcase
casez ({new_n151_, new_n509_, new_n2703_})
3'b11? : new_n4131_ = 1'b1;
3'b??1 : new_n4131_ = 1'b1;
default : new_n4131_ = 1'b0;
endcase
casez ({new_n1027_, new_n2704_})
2'b00 : new_n4132_ = 1'b1;
default : new_n4132_ = 1'b0;
endcase
casez ({new_n606_, new_n634_})
2'b00 : new_n4133_ = 1'b1;
default : new_n4133_ = 1'b0;
endcase
casez ({new_n676_, new_n2707_})
2'b00 : new_n4134_ = 1'b1;
default : new_n4134_ = 1'b0;
endcase
casez ({new_n137_, new_n401_, new_n2708_})
3'b11? : new_n4135_ = 1'b1;
3'b??1 : new_n4135_ = 1'b1;
default : new_n4135_ = 1'b0;
endcase
casez ({new_n1593_, new_n2709_})
2'b00 : new_n4136_ = 1'b1;
default : new_n4136_ = 1'b0;
endcase
casez ({new_n2571_, new_n2710_})
2'b00 : new_n4137_ = 1'b1;
default : new_n4137_ = 1'b0;
endcase
casez ({new_n861_, new_n2710_})
2'b00 : new_n4138_ = 1'b1;
default : new_n4138_ = 1'b0;
endcase
casez ({new_n107_, new_n215_, new_n635_})
3'b01? : new_n4139_ = 1'b1;
3'b??1 : new_n4139_ = 1'b1;
default : new_n4139_ = 1'b0;
endcase
casez ({new_n1638_, new_n2714_})
2'b00 : new_n4140_ = 1'b1;
default : new_n4140_ = 1'b0;
endcase
casez ({new_n187_, new_n961_, new_n199_, new_n2716_})
4'b11?? : new_n4141_ = 1'b1;
4'b??11 : new_n4141_ = 1'b1;
default : new_n4141_ = 1'b0;
endcase
casez ({new_n1036_, new_n2717_})
2'b00 : new_n4142_ = 1'b1;
default : new_n4142_ = 1'b0;
endcase
casez ({new_n112_, new_n301_, new_n2717_})
3'b11? : new_n4143_ = 1'b1;
3'b??1 : new_n4143_ = 1'b1;
default : new_n4143_ = 1'b0;
endcase
casez ({new_n177_, new_n207_, new_n2718_})
3'b11? : new_n4144_ = 1'b1;
3'b??1 : new_n4144_ = 1'b1;
default : new_n4144_ = 1'b0;
endcase
casez ({new_n945_, new_n2719_})
2'b00 : new_n4145_ = 1'b1;
default : new_n4145_ = 1'b0;
endcase
casez ({new_n2653_, new_n2719_})
2'b00 : new_n4146_ = 1'b1;
default : new_n4146_ = 1'b0;
endcase
casez ({new_n179_, new_n417_, new_n2720_})
3'b11? : new_n4147_ = 1'b1;
3'b??1 : new_n4147_ = 1'b1;
default : new_n4147_ = 1'b0;
endcase
casez ({new_n230_, new_n428_, new_n2723_})
3'b10? : new_n4148_ = 1'b1;
3'b??1 : new_n4148_ = 1'b1;
default : new_n4148_ = 1'b0;
endcase
casez ({new_n1899_, new_n2724_})
2'b00 : new_n4149_ = 1'b1;
default : new_n4149_ = 1'b0;
endcase
casez ({new_n4650_, new_n636_})
2'b1? : new_n4150_ = 1'b1;
2'b?1 : new_n4150_ = 1'b1;
default : new_n4150_ = 1'b0;
endcase
casez ({new_n1364_, new_n2725_})
2'b00 : new_n4151_ = 1'b1;
default : new_n4151_ = 1'b0;
endcase
casez ({new_n869_, new_n2726_})
2'b00 : new_n4152_ = 1'b1;
default : new_n4152_ = 1'b0;
endcase
casez ({new_n1151_, new_n2727_})
2'b00 : new_n4153_ = 1'b1;
default : new_n4153_ = 1'b0;
endcase
casez ({new_n784_, new_n2728_})
2'b00 : new_n4154_ = 1'b1;
default : new_n4154_ = 1'b0;
endcase
casez ({new_n1852_, new_n2728_})
2'b00 : new_n4155_ = 1'b1;
default : new_n4155_ = 1'b0;
endcase
casez ({new_n230_, new_n356_, new_n2730_})
3'b11? : new_n4156_ = 1'b1;
3'b??1 : new_n4156_ = 1'b1;
default : new_n4156_ = 1'b0;
endcase
casez ({new_n150_, new_n465_, new_n2731_})
3'b10? : new_n4157_ = 1'b1;
3'b??1 : new_n4157_ = 1'b1;
default : new_n4157_ = 1'b0;
endcase
casez ({new_n1115_, new_n2734_})
2'b00 : new_n4158_ = 1'b1;
default : new_n4158_ = 1'b0;
endcase
casez ({new_n1612_, new_n2735_})
2'b00 : new_n4159_ = 1'b1;
default : new_n4159_ = 1'b0;
endcase
casez ({new_n245_, new_n955_})
2'b00 : new_n4160_ = 1'b1;
default : new_n4160_ = 1'b0;
endcase
casez ({new_n4662_, new_n638_})
2'b1? : new_n4161_ = 1'b1;
2'b?1 : new_n4161_ = 1'b1;
default : new_n4161_ = 1'b0;
endcase
casez ({new_n1829_, new_n2738_})
2'b00 : new_n4162_ = 1'b1;
default : new_n4162_ = 1'b0;
endcase
casez ({new_n139_, new_n2739_})
2'b00 : new_n4163_ = 1'b1;
default : new_n4163_ = 1'b0;
endcase
casez ({new_n391_, new_n2742_})
2'b00 : new_n4164_ = 1'b1;
default : new_n4164_ = 1'b0;
endcase
casez ({new_n1960_, new_n2743_})
2'b00 : new_n4165_ = 1'b1;
default : new_n4165_ = 1'b0;
endcase
casez ({new_n1043_, new_n2744_})
2'b00 : new_n4166_ = 1'b1;
default : new_n4166_ = 1'b0;
endcase
casez ({new_n1588_, new_n2744_})
2'b00 : new_n4167_ = 1'b1;
default : new_n4167_ = 1'b0;
endcase
casez ({new_n223_, new_n508_, new_n2745_})
3'b11? : new_n4168_ = 1'b1;
3'b??1 : new_n4168_ = 1'b1;
default : new_n4168_ = 1'b0;
endcase
casez ({new_n740_, new_n2746_})
2'b00 : new_n4169_ = 1'b1;
default : new_n4169_ = 1'b0;
endcase
casez ({new_n89_, new_n162_, new_n2751_})
3'b11? : new_n4170_ = 1'b1;
3'b??1 : new_n4170_ = 1'b1;
default : new_n4170_ = 1'b0;
endcase
casez ({x[0], new_n958_, new_n142_, new_n302_})
4'b11?? : new_n4171_ = 1'b1;
4'b??10 : new_n4171_ = 1'b1;
default : new_n4171_ = 1'b0;
endcase
casez ({new_n2639_, new_n2752_})
2'b00 : new_n4172_ = 1'b1;
default : new_n4172_ = 1'b0;
endcase
casez ({new_n223_, new_n257_, new_n2752_})
3'b11? : new_n4173_ = 1'b1;
3'b??1 : new_n4173_ = 1'b1;
default : new_n4173_ = 1'b0;
endcase
casez ({new_n4610_, new_n959_})
2'b1? : new_n4174_ = 1'b1;
2'b?1 : new_n4174_ = 1'b1;
default : new_n4174_ = 1'b0;
endcase
casez ({new_n335_, new_n2755_})
2'b00 : new_n4175_ = 1'b1;
default : new_n4175_ = 1'b0;
endcase
casez ({new_n335_, new_n2756_})
2'b00 : new_n4176_ = 1'b1;
default : new_n4176_ = 1'b0;
endcase
casez ({new_n86_, new_n1159_, new_n2758_})
3'b11? : new_n4177_ = 1'b1;
3'b??1 : new_n4177_ = 1'b1;
default : new_n4177_ = 1'b0;
endcase
casez ({new_n717_, new_n959_})
2'b00 : new_n4178_ = 1'b1;
default : new_n4178_ = 1'b0;
endcase
casez ({new_n451_, new_n639_})
2'b00 : new_n4179_ = 1'b1;
default : new_n4179_ = 1'b0;
endcase
casez ({new_n1846_, new_n2761_})
2'b00 : new_n4180_ = 1'b1;
default : new_n4180_ = 1'b0;
endcase
casez ({new_n1638_, new_n2763_})
2'b00 : new_n4181_ = 1'b1;
default : new_n4181_ = 1'b0;
endcase
casez ({new_n424_, new_n2765_})
2'b00 : new_n4182_ = 1'b1;
default : new_n4182_ = 1'b0;
endcase
casez ({new_n2761_, new_n2766_})
2'b00 : new_n4183_ = 1'b1;
default : new_n4183_ = 1'b0;
endcase
casez ({y[2], new_n491_, new_n960_})
3'b10? : new_n4184_ = 1'b1;
3'b??1 : new_n4184_ = 1'b1;
default : new_n4184_ = 1'b0;
endcase
casez ({new_n301_, new_n961_, new_n308_, new_n321_})
4'b11?? : new_n4185_ = 1'b1;
4'b??11 : new_n4185_ = 1'b1;
default : new_n4185_ = 1'b0;
endcase
casez ({new_n340_, new_n2769_})
2'b00 : new_n4186_ = 1'b1;
default : new_n4186_ = 1'b0;
endcase
casez ({new_n743_, new_n962_})
2'b00 : new_n4187_ = 1'b1;
default : new_n4187_ = 1'b0;
endcase
casez ({new_n118_, new_n2538_, new_n2772_})
3'b10? : new_n4188_ = 1'b1;
3'b??1 : new_n4188_ = 1'b1;
default : new_n4188_ = 1'b0;
endcase
casez ({new_n1607_, new_n2776_})
2'b00 : new_n4189_ = 1'b1;
default : new_n4189_ = 1'b0;
endcase
casez ({new_n1130_, new_n2776_})
2'b00 : new_n4190_ = 1'b1;
default : new_n4190_ = 1'b0;
endcase
casez ({new_n858_, new_n963_})
2'b00 : new_n4191_ = 1'b1;
default : new_n4191_ = 1'b0;
endcase
casez ({new_n83_, new_n104_, new_n963_})
3'b11? : new_n4192_ = 1'b1;
3'b??1 : new_n4192_ = 1'b1;
default : new_n4192_ = 1'b0;
endcase
casez ({new_n1046_, new_n2779_})
2'b00 : new_n4193_ = 1'b1;
default : new_n4193_ = 1'b0;
endcase
casez ({new_n620_, new_n2779_})
2'b00 : new_n4194_ = 1'b1;
default : new_n4194_ = 1'b0;
endcase
casez ({new_n187_, new_n444_, new_n963_})
3'b11? : new_n4195_ = 1'b1;
3'b??1 : new_n4195_ = 1'b1;
default : new_n4195_ = 1'b0;
endcase
casez ({new_n382_, new_n963_})
2'b00 : new_n4196_ = 1'b1;
default : new_n4196_ = 1'b0;
endcase
casez ({new_n536_, new_n964_})
2'b00 : new_n4197_ = 1'b1;
default : new_n4197_ = 1'b0;
endcase
casez ({new_n88_, new_n155_, new_n353_})
3'b11? : new_n4198_ = 1'b1;
3'b??1 : new_n4198_ = 1'b1;
default : new_n4198_ = 1'b0;
endcase
casez ({new_n132_, new_n201_, new_n157_, new_n200_})
4'b11?? : new_n4199_ = 1'b1;
4'b??11 : new_n4199_ = 1'b1;
default : new_n4199_ = 1'b0;
endcase
casez ({new_n244_, new_n364_})
2'b01 : new_n4200_ = 1'b1;
default : new_n4200_ = 1'b0;
endcase
casez ({new_n525_, new_n1542_})
2'b00 : new_n4201_ = 1'b1;
default : new_n4201_ = 1'b0;
endcase
casez ({new_n1134_, new_n1542_})
2'b00 : new_n4202_ = 1'b1;
default : new_n4202_ = 1'b0;
endcase
casez ({new_n414_, new_n1543_})
2'b00 : new_n4203_ = 1'b1;
default : new_n4203_ = 1'b0;
endcase
casez ({new_n871_, new_n1543_})
2'b00 : new_n4204_ = 1'b1;
default : new_n4204_ = 1'b0;
endcase
casez ({new_n677_, new_n728_, new_n1544_})
3'b1?? : new_n4205_ = 1'b1;
3'b?11 : new_n4205_ = 1'b1;
default : new_n4205_ = 1'b0;
endcase
casez ({new_n243_, new_n1545_, new_n1121_})
3'b11? : new_n4206_ = 1'b1;
3'b??1 : new_n4206_ = 1'b1;
default : new_n4206_ = 1'b0;
endcase
casez ({new_n162_, new_n1303_, new_n321_, new_n1552_})
4'b10?? : new_n4207_ = 1'b1;
4'b??10 : new_n4207_ = 1'b1;
default : new_n4207_ = 1'b0;
endcase
casez ({new_n99_, new_n356_, new_n1554_})
3'b01? : new_n4208_ = 1'b1;
3'b??0 : new_n4208_ = 1'b1;
default : new_n4208_ = 1'b0;
endcase
casez ({new_n156_, new_n1557_})
2'b00 : new_n4209_ = 1'b1;
default : new_n4209_ = 1'b0;
endcase
casez ({new_n963_, new_n1557_})
2'b00 : new_n4210_ = 1'b1;
default : new_n4210_ = 1'b0;
endcase
casez ({new_n438_, new_n2924_})
2'b00 : new_n4211_ = 1'b1;
default : new_n4211_ = 1'b0;
endcase
casez ({new_n2583_, new_n2940_})
2'b00 : new_n4212_ = 1'b1;
default : new_n4212_ = 1'b0;
endcase
casez ({new_n1645_, new_n2942_})
2'b00 : new_n4213_ = 1'b1;
default : new_n4213_ = 1'b0;
endcase
casez ({new_n675_, new_n2943_})
2'b00 : new_n4214_ = 1'b1;
default : new_n4214_ = 1'b0;
endcase
casez ({new_n716_, new_n2947_})
2'b00 : new_n4215_ = 1'b1;
default : new_n4215_ = 1'b0;
endcase
casez ({new_n1342_, new_n2953_})
2'b00 : new_n4216_ = 1'b1;
default : new_n4216_ = 1'b0;
endcase
casez ({new_n104_, new_n250_, new_n1563_})
3'b11? : new_n4217_ = 1'b1;
3'b??1 : new_n4217_ = 1'b1;
default : new_n4217_ = 1'b0;
endcase
casez ({new_n751_, new_n2956_})
2'b00 : new_n4218_ = 1'b1;
default : new_n4218_ = 1'b0;
endcase
casez ({new_n414_, new_n2957_})
2'b00 : new_n4219_ = 1'b1;
default : new_n4219_ = 1'b0;
endcase
casez ({new_n305_, new_n417_, new_n1563_})
3'b11? : new_n4220_ = 1'b1;
3'b??1 : new_n4220_ = 1'b1;
default : new_n4220_ = 1'b0;
endcase
casez ({new_n620_, new_n1564_})
2'b00 : new_n4221_ = 1'b1;
default : new_n4221_ = 1'b0;
endcase
casez ({new_n742_, new_n2965_})
2'b00 : new_n4222_ = 1'b1;
default : new_n4222_ = 1'b0;
endcase
casez ({new_n310_, new_n2965_})
2'b00 : new_n4223_ = 1'b1;
default : new_n4223_ = 1'b0;
endcase
casez ({new_n1172_, new_n2970_})
2'b00 : new_n4224_ = 1'b1;
default : new_n4224_ = 1'b0;
endcase
casez ({new_n752_, new_n2972_})
2'b00 : new_n4225_ = 1'b1;
default : new_n4225_ = 1'b0;
endcase
casez ({new_n87_, new_n2975_, new_n2775_})
3'b11? : new_n4226_ = 1'b1;
3'b??1 : new_n4226_ = 1'b1;
default : new_n4226_ = 1'b0;
endcase
casez ({new_n325_, new_n668_})
2'b00 : new_n4227_ = 1'b1;
default : new_n4227_ = 1'b0;
endcase
casez ({new_n1162_, new_n2979_})
2'b00 : new_n4228_ = 1'b1;
default : new_n4228_ = 1'b0;
endcase
casez ({new_n81_, new_n1175_, new_n102_, new_n2980_})
4'b01?? : new_n4229_ = 1'b1;
4'b??11 : new_n4229_ = 1'b1;
default : new_n4229_ = 1'b0;
endcase
casez ({new_n676_, new_n1568_})
2'b00 : new_n4230_ = 1'b1;
default : new_n4230_ = 1'b0;
endcase
casez ({new_n1264_, new_n2986_})
2'b01 : new_n4231_ = 1'b1;
default : new_n4231_ = 1'b0;
endcase
casez ({new_n535_, new_n668_})
2'b00 : new_n4232_ = 1'b1;
default : new_n4232_ = 1'b0;
endcase
casez ({new_n79_, new_n97_, new_n222_, new_n1569_})
4'b101? : new_n4233_ = 1'b1;
4'b???1 : new_n4233_ = 1'b1;
default : new_n4233_ = 1'b0;
endcase
casez ({new_n179_, new_n1570_, new_n784_})
3'b11? : new_n4234_ = 1'b1;
3'b??1 : new_n4234_ = 1'b1;
default : new_n4234_ = 1'b0;
endcase
casez ({new_n487_, new_n999_})
2'b01 : new_n4235_ = 1'b1;
default : new_n4235_ = 1'b0;
endcase
casez ({new_n4652_, new_n338_, new_n370_})
3'b1?? : new_n4236_ = 1'b1;
3'b?10 : new_n4236_ = 1'b1;
default : new_n4236_ = 1'b0;
endcase
casez ({new_n311_, new_n1002_})
2'b00 : new_n4237_ = 1'b1;
default : new_n4237_ = 1'b0;
endcase
casez ({new_n1358_, new_n1571_})
2'b00 : new_n4238_ = 1'b1;
default : new_n4238_ = 1'b0;
endcase
casez ({new_n683_, new_n1002_})
2'b00 : new_n4239_ = 1'b1;
default : new_n4239_ = 1'b0;
endcase
casez ({new_n184_, new_n214_, new_n1003_})
3'b11? : new_n4240_ = 1'b1;
3'b??1 : new_n4240_ = 1'b1;
default : new_n4240_ = 1'b0;
endcase
casez ({new_n1118_, new_n1572_})
2'b00 : new_n4241_ = 1'b1;
default : new_n4241_ = 1'b0;
endcase
casez ({new_n231_, new_n3017_})
2'b01 : new_n4242_ = 1'b1;
default : new_n4242_ = 1'b0;
endcase
casez ({new_n540_, new_n1573_})
2'b00 : new_n4243_ = 1'b1;
default : new_n4243_ = 1'b0;
endcase
casez ({new_n858_, new_n1573_})
2'b00 : new_n4244_ = 1'b1;
default : new_n4244_ = 1'b0;
endcase
casez ({new_n854_, new_n1574_})
2'b00 : new_n4245_ = 1'b1;
default : new_n4245_ = 1'b0;
endcase
casez ({new_n1105_, new_n1574_})
2'b00 : new_n4246_ = 1'b1;
default : new_n4246_ = 1'b0;
endcase
casez ({new_n190_, new_n216_, new_n1574_})
3'b11? : new_n4247_ = 1'b1;
3'b??1 : new_n4247_ = 1'b1;
default : new_n4247_ = 1'b0;
endcase
casez ({v[1], new_n1005_, new_n209_, new_n421_})
4'b01?? : new_n4248_ = 1'b1;
4'b??11 : new_n4248_ = 1'b1;
default : new_n4248_ = 1'b0;
endcase
casez ({new_n939_, new_n1576_})
2'b00 : new_n4249_ = 1'b1;
default : new_n4249_ = 1'b0;
endcase
casez ({new_n482_, new_n1007_})
2'b00 : new_n4250_ = 1'b1;
default : new_n4250_ = 1'b0;
endcase
casez ({y[2], new_n927_, new_n3054_})
3'b11? : new_n4251_ = 1'b1;
3'b??0 : new_n4251_ = 1'b1;
default : new_n4251_ = 1'b0;
endcase
casez ({new_n115_, new_n123_, new_n1007_})
3'b11? : new_n4252_ = 1'b1;
3'b??1 : new_n4252_ = 1'b1;
default : new_n4252_ = 1'b0;
endcase
casez ({new_n250_, new_n1159_, new_n321_, new_n1580_})
4'b11?? : new_n4253_ = 1'b1;
4'b??11 : new_n4253_ = 1'b1;
default : new_n4253_ = 1'b0;
endcase
casez ({new_n177_, new_n264_, new_n1009_})
3'b11? : new_n4254_ = 1'b1;
3'b??1 : new_n4254_ = 1'b1;
default : new_n4254_ = 1'b0;
endcase
casez ({new_n79_, new_n189_, new_n1582_})
3'b11? : new_n4255_ = 1'b1;
3'b??1 : new_n4255_ = 1'b1;
default : new_n4255_ = 1'b0;
endcase
casez ({new_n602_, new_n675_})
2'b00 : new_n4256_ = 1'b1;
default : new_n4256_ = 1'b0;
endcase
casez ({new_n1105_, new_n1582_})
2'b00 : new_n4257_ = 1'b1;
default : new_n4257_ = 1'b0;
endcase
casez ({new_n387_, new_n1583_})
2'b00 : new_n4258_ = 1'b1;
default : new_n4258_ = 1'b0;
endcase
casez ({new_n290_, new_n1583_})
2'b00 : new_n4259_ = 1'b1;
default : new_n4259_ = 1'b0;
endcase
casez ({new_n101_, new_n244_, new_n377_})
3'b11? : new_n4260_ = 1'b1;
3'b??1 : new_n4260_ = 1'b1;
default : new_n4260_ = 1'b0;
endcase
casez ({new_n1004_, new_n1584_})
2'b00 : new_n4261_ = 1'b1;
default : new_n4261_ = 1'b0;
endcase
casez ({new_n208_, new_n369_, new_n1010_})
3'b11? : new_n4262_ = 1'b1;
3'b??1 : new_n4262_ = 1'b1;
default : new_n4262_ = 1'b0;
endcase
casez ({new_n139_, new_n307_, new_n1584_})
3'b11? : new_n4263_ = 1'b1;
3'b??1 : new_n4263_ = 1'b1;
default : new_n4263_ = 1'b0;
endcase
casez ({x[0], new_n527_, new_n1586_})
3'b01? : new_n4264_ = 1'b1;
3'b??1 : new_n4264_ = 1'b1;
default : new_n4264_ = 1'b0;
endcase
casez ({new_n4637_, new_n1587_})
2'b1? : new_n4265_ = 1'b1;
2'b?1 : new_n4265_ = 1'b1;
default : new_n4265_ = 1'b0;
endcase
casez ({new_n115_, new_n240_, new_n1011_})
3'b11? : new_n4266_ = 1'b1;
3'b??1 : new_n4266_ = 1'b1;
default : new_n4266_ = 1'b0;
endcase
casez ({new_n1136_, new_n1588_})
2'b00 : new_n4267_ = 1'b1;
default : new_n4267_ = 1'b0;
endcase
casez ({new_n4591_, new_n1588_})
2'b1? : new_n4268_ = 1'b1;
2'b?1 : new_n4268_ = 1'b1;
default : new_n4268_ = 1'b0;
endcase
casez ({new_n4654_, new_n325_})
2'b1? : new_n4269_ = 1'b1;
2'b?1 : new_n4269_ = 1'b1;
default : new_n4269_ = 1'b0;
endcase
casez ({new_n208_, new_n398_, new_n677_})
3'b11? : new_n4270_ = 1'b1;
3'b??1 : new_n4270_ = 1'b1;
default : new_n4270_ = 1'b0;
endcase
casez ({new_n790_, new_n1589_})
2'b00 : new_n4271_ = 1'b1;
default : new_n4271_ = 1'b0;
endcase
casez ({new_n471_, new_n1012_})
2'b00 : new_n4272_ = 1'b1;
default : new_n4272_ = 1'b0;
endcase
casez ({u[1], new_n1013_, new_n85_, new_n606_})
4'b01?? : new_n4273_ = 1'b1;
4'b??11 : new_n4273_ = 1'b1;
default : new_n4273_ = 1'b0;
endcase
casez ({new_n137_, new_n381_})
2'b00 : new_n4274_ = 1'b1;
default : new_n4274_ = 1'b0;
endcase
casez ({new_n4612_, new_n1014_})
2'b1? : new_n4275_ = 1'b1;
2'b?1 : new_n4275_ = 1'b1;
default : new_n4275_ = 1'b0;
endcase
casez ({new_n229_, new_n287_, new_n1591_})
3'b11? : new_n4276_ = 1'b1;
3'b??1 : new_n4276_ = 1'b1;
default : new_n4276_ = 1'b0;
endcase
casez ({new_n947_, new_n1014_})
2'b00 : new_n4277_ = 1'b1;
default : new_n4277_ = 1'b0;
endcase
casez ({new_n780_, new_n1593_})
2'b00 : new_n4278_ = 1'b1;
default : new_n4278_ = 1'b0;
endcase
casez ({new_n941_, new_n1595_})
2'b00 : new_n4279_ = 1'b1;
default : new_n4279_ = 1'b0;
endcase
casez ({new_n639_, new_n1595_})
2'b00 : new_n4280_ = 1'b1;
default : new_n4280_ = 1'b0;
endcase
casez ({new_n584_, new_n679_})
2'b00 : new_n4281_ = 1'b1;
default : new_n4281_ = 1'b0;
endcase
casez ({x[2], new_n114_, new_n1016_})
3'b11? : new_n4282_ = 1'b1;
3'b??1 : new_n4282_ = 1'b1;
default : new_n4282_ = 1'b0;
endcase
casez ({new_n1027_, new_n1596_})
2'b00 : new_n4283_ = 1'b1;
default : new_n4283_ = 1'b0;
endcase
casez ({new_n122_, new_n213_})
2'b00 : new_n4284_ = 1'b1;
default : new_n4284_ = 1'b0;
endcase
casez ({new_n454_, new_n1016_})
2'b00 : new_n4285_ = 1'b1;
default : new_n4285_ = 1'b0;
endcase
casez ({new_n1140_, new_n1598_})
2'b00 : new_n4286_ = 1'b1;
default : new_n4286_ = 1'b0;
endcase
casez ({new_n220_, new_n469_, new_n1598_})
3'b11? : new_n4287_ = 1'b1;
3'b??1 : new_n4287_ = 1'b1;
default : new_n4287_ = 1'b0;
endcase
casez ({new_n460_, new_n680_})
2'b00 : new_n4288_ = 1'b1;
default : new_n4288_ = 1'b0;
endcase
casez ({new_n414_, new_n3210_})
2'b01 : new_n4289_ = 1'b1;
default : new_n4289_ = 1'b0;
endcase
casez ({new_n1124_, new_n1599_})
2'b00 : new_n4290_ = 1'b1;
default : new_n4290_ = 1'b0;
endcase
casez ({new_n192_, new_n1100_, new_n1600_})
3'b10? : new_n4291_ = 1'b1;
3'b??1 : new_n4291_ = 1'b1;
default : new_n4291_ = 1'b0;
endcase
casez ({new_n89_, new_n435_, new_n1601_})
3'b11? : new_n4292_ = 1'b1;
3'b??1 : new_n4292_ = 1'b1;
default : new_n4292_ = 1'b0;
endcase
casez ({new_n552_, new_n682_})
2'b00 : new_n4293_ = 1'b1;
default : new_n4293_ = 1'b0;
endcase
casez ({new_n1009_, new_n1602_})
2'b00 : new_n4294_ = 1'b1;
default : new_n4294_ = 1'b0;
endcase
casez ({new_n668_, new_n1018_})
2'b00 : new_n4295_ = 1'b1;
default : new_n4295_ = 1'b0;
endcase
casez ({new_n472_, new_n1603_})
2'b00 : new_n4296_ = 1'b1;
default : new_n4296_ = 1'b0;
endcase
casez ({new_n1012_, new_n1603_})
2'b00 : new_n4297_ = 1'b1;
default : new_n4297_ = 1'b0;
endcase
casez ({new_n859_, new_n1604_})
2'b00 : new_n4298_ = 1'b1;
default : new_n4298_ = 1'b0;
endcase
casez ({new_n540_, new_n1604_})
2'b00 : new_n4299_ = 1'b1;
default : new_n4299_ = 1'b0;
endcase
casez ({new_n543_, new_n1606_})
2'b00 : new_n4300_ = 1'b1;
default : new_n4300_ = 1'b0;
endcase
casez ({new_n1365_, new_n1606_})
2'b00 : new_n4301_ = 1'b1;
default : new_n4301_ = 1'b0;
endcase
casez ({new_n603_, new_n1021_})
2'b00 : new_n4302_ = 1'b1;
default : new_n4302_ = 1'b0;
endcase
casez ({new_n442_, new_n683_})
2'b00 : new_n4303_ = 1'b1;
default : new_n4303_ = 1'b0;
endcase
casez ({new_n162_, new_n210_, new_n1022_})
3'b11? : new_n4304_ = 1'b1;
3'b??1 : new_n4304_ = 1'b1;
default : new_n4304_ = 1'b0;
endcase
casez ({new_n1097_, new_n3284_})
2'b01 : new_n4305_ = 1'b1;
default : new_n4305_ = 1'b0;
endcase
casez ({new_n4615_, new_n330_})
2'b1? : new_n4306_ = 1'b1;
2'b?1 : new_n4306_ = 1'b1;
default : new_n4306_ = 1'b0;
endcase
casez ({new_n737_, new_n1022_})
2'b00 : new_n4307_ = 1'b1;
default : new_n4307_ = 1'b0;
endcase
casez ({new_n88_, new_n340_, new_n1022_})
3'b01? : new_n4308_ = 1'b1;
3'b??1 : new_n4308_ = 1'b1;
default : new_n4308_ = 1'b0;
endcase
casez ({new_n1179_, new_n1610_})
2'b00 : new_n4309_ = 1'b1;
default : new_n4309_ = 1'b0;
endcase
casez ({new_n584_, new_n1023_})
2'b00 : new_n4310_ = 1'b1;
default : new_n4310_ = 1'b0;
endcase
casez ({new_n139_, new_n319_, new_n1611_})
3'b10? : new_n4311_ = 1'b1;
3'b??1 : new_n4311_ = 1'b1;
default : new_n4311_ = 1'b0;
endcase
casez ({new_n88_, new_n1024_, new_n146_, new_n156_})
4'b11?? : new_n4312_ = 1'b1;
4'b??11 : new_n4312_ = 1'b1;
default : new_n4312_ = 1'b0;
endcase
casez ({new_n86_, new_n1025_, new_n944_})
3'b01? : new_n4313_ = 1'b1;
3'b??1 : new_n4313_ = 1'b1;
default : new_n4313_ = 1'b0;
endcase
casez ({new_n249_, new_n388_})
2'b00 : new_n4314_ = 1'b1;
default : new_n4314_ = 1'b0;
endcase
casez ({x[0], new_n669_, new_n1026_})
3'b01? : new_n4315_ = 1'b1;
3'b??1 : new_n4315_ = 1'b1;
default : new_n4315_ = 1'b0;
endcase
casez ({new_n2591_, new_n3324_})
2'b00 : new_n4316_ = 1'b1;
default : new_n4316_ = 1'b0;
endcase
casez ({new_n1115_, new_n1616_})
2'b00 : new_n4317_ = 1'b1;
default : new_n4317_ = 1'b0;
endcase
casez ({v[1], new_n1396_, new_n3325_})
3'b11? : new_n4318_ = 1'b1;
3'b??1 : new_n4318_ = 1'b1;
default : new_n4318_ = 1'b0;
endcase
casez ({new_n1009_, new_n1027_})
2'b00 : new_n4319_ = 1'b1;
default : new_n4319_ = 1'b0;
endcase
casez ({new_n1141_, new_n3328_})
2'b00 : new_n4320_ = 1'b1;
default : new_n4320_ = 1'b0;
endcase
casez ({new_n2638_, new_n3331_})
2'b00 : new_n4321_ = 1'b1;
default : new_n4321_ = 1'b0;
endcase
casez ({new_n1144_, new_n3331_})
2'b00 : new_n4322_ = 1'b1;
default : new_n4322_ = 1'b0;
endcase
casez ({new_n4617_, new_n224_, new_n243_})
3'b1?? : new_n4323_ = 1'b1;
3'b?11 : new_n4323_ = 1'b1;
default : new_n4323_ = 1'b0;
endcase
casez ({new_n1017_, new_n3337_})
2'b00 : new_n4324_ = 1'b1;
default : new_n4324_ = 1'b0;
endcase
casez ({v[1], new_n602_, new_n1028_})
3'b01? : new_n4325_ = 1'b1;
3'b??1 : new_n4325_ = 1'b1;
default : new_n4325_ = 1'b0;
endcase
casez ({new_n1894_, new_n3339_})
2'b00 : new_n4326_ = 1'b1;
default : new_n4326_ = 1'b0;
endcase
casez ({new_n1346_, new_n1618_})
2'b00 : new_n4327_ = 1'b1;
default : new_n4327_ = 1'b0;
endcase
casez ({new_n1612_, new_n3340_})
2'b00 : new_n4328_ = 1'b1;
default : new_n4328_ = 1'b0;
endcase
casez ({new_n1260_, new_n1619_})
2'b00 : new_n4329_ = 1'b1;
default : new_n4329_ = 1'b0;
endcase
casez ({new_n1132_, new_n3342_})
2'b00 : new_n4330_ = 1'b1;
default : new_n4330_ = 1'b0;
endcase
casez ({v[1], new_n234_, new_n101_, new_n1620_})
4'b11?? : new_n4331_ = 1'b1;
4'b??11 : new_n4331_ = 1'b1;
default : new_n4331_ = 1'b0;
endcase
casez ({new_n1833_, new_n3344_})
2'b00 : new_n4332_ = 1'b1;
default : new_n4332_ = 1'b0;
endcase
casez ({new_n1853_, new_n3345_})
2'b00 : new_n4333_ = 1'b1;
default : new_n4333_ = 1'b0;
endcase
casez ({new_n345_, new_n1029_})
2'b00 : new_n4334_ = 1'b1;
default : new_n4334_ = 1'b0;
endcase
casez ({new_n267_, new_n3347_, new_n422_, new_n441_})
4'b11?? : new_n4335_ = 1'b1;
4'b??11 : new_n4335_ = 1'b1;
default : new_n4335_ = 1'b0;
endcase
casez ({y[1], new_n619_, new_n318_, new_n1620_})
4'b11?? : new_n4336_ = 1'b1;
4'b??11 : new_n4336_ = 1'b1;
default : new_n4336_ = 1'b0;
endcase
casez ({new_n85_, new_n139_, new_n1029_})
3'b01? : new_n4337_ = 1'b1;
3'b??1 : new_n4337_ = 1'b1;
default : new_n4337_ = 1'b0;
endcase
casez ({new_n553_, new_n1030_})
2'b00 : new_n4338_ = 1'b1;
default : new_n4338_ = 1'b0;
endcase
casez ({new_n1836_, new_n3351_})
2'b00 : new_n4339_ = 1'b1;
default : new_n4339_ = 1'b0;
endcase
casez ({new_n1597_, new_n3351_})
2'b00 : new_n4340_ = 1'b1;
default : new_n4340_ = 1'b0;
endcase
casez ({new_n361_, new_n391_})
2'b00 : new_n4341_ = 1'b1;
default : new_n4341_ = 1'b0;
endcase
casez ({new_n1111_, new_n3355_})
2'b00 : new_n4342_ = 1'b1;
default : new_n4342_ = 1'b0;
endcase
casez ({new_n240_, new_n273_, new_n1030_})
3'b11? : new_n4343_ = 1'b1;
3'b??1 : new_n4343_ = 1'b1;
default : new_n4343_ = 1'b0;
endcase
casez ({new_n784_, new_n3358_})
2'b00 : new_n4344_ = 1'b1;
default : new_n4344_ = 1'b0;
endcase
casez ({new_n1841_, new_n3362_})
2'b00 : new_n4345_ = 1'b1;
default : new_n4345_ = 1'b0;
endcase
casez ({new_n855_, new_n3364_})
2'b00 : new_n4346_ = 1'b1;
default : new_n4346_ = 1'b0;
endcase
casez ({new_n1044_, new_n1623_})
2'b00 : new_n4347_ = 1'b1;
default : new_n4347_ = 1'b0;
endcase
casez ({new_n4627_, new_n3365_})
2'b1? : new_n4348_ = 1'b1;
2'b?1 : new_n4348_ = 1'b1;
default : new_n4348_ = 1'b0;
endcase
casez ({new_n245_, new_n1031_})
2'b00 : new_n4349_ = 1'b1;
default : new_n4349_ = 1'b0;
endcase
casez ({new_n2746_, new_n3369_})
2'b00 : new_n4350_ = 1'b1;
default : new_n4350_ = 1'b0;
endcase
casez ({new_n83_, new_n2689_, new_n3371_})
3'b11? : new_n4351_ = 1'b1;
3'b??1 : new_n4351_ = 1'b1;
default : new_n4351_ = 1'b0;
endcase
casez ({new_n2633_, new_n3374_})
2'b00 : new_n4352_ = 1'b1;
default : new_n4352_ = 1'b0;
endcase
casez ({new_n282_, new_n3375_})
2'b00 : new_n4353_ = 1'b1;
default : new_n4353_ = 1'b0;
endcase
casez ({new_n2591_, new_n3379_})
2'b00 : new_n4354_ = 1'b1;
default : new_n4354_ = 1'b0;
endcase
casez ({new_n583_, new_n3382_})
2'b00 : new_n4355_ = 1'b1;
default : new_n4355_ = 1'b0;
endcase
casez ({new_n1945_, new_n3383_})
2'b00 : new_n4356_ = 1'b1;
default : new_n4356_ = 1'b0;
endcase
casez ({v[0], new_n105_, new_n3384_})
3'b11? : new_n4357_ = 1'b1;
3'b??1 : new_n4357_ = 1'b1;
default : new_n4357_ = 1'b0;
endcase
casez ({new_n122_, new_n217_})
2'b00 : new_n4358_ = 1'b1;
default : new_n4358_ = 1'b0;
endcase
casez ({new_n747_, new_n1626_})
2'b00 : new_n4359_ = 1'b1;
default : new_n4359_ = 1'b0;
endcase
casez ({x[0], new_n3387_, new_n150_, new_n372_})
4'b11?? : new_n4360_ = 1'b1;
4'b??11 : new_n4360_ = 1'b1;
default : new_n4360_ = 1'b0;
endcase
casez ({new_n396_, new_n1626_})
2'b00 : new_n4361_ = 1'b1;
default : new_n4361_ = 1'b0;
endcase
casez ({new_n1139_, new_n1627_})
2'b00 : new_n4362_ = 1'b1;
default : new_n4362_ = 1'b0;
endcase
casez ({new_n1862_, new_n3396_})
2'b00 : new_n4363_ = 1'b1;
default : new_n4363_ = 1'b0;
endcase
casez ({new_n2652_, new_n3398_, new_n2932_, new_n3389_})
4'b11?? : new_n4364_ = 1'b1;
4'b??11 : new_n4364_ = 1'b1;
default : new_n4364_ = 1'b0;
endcase
casez ({new_n1017_, new_n3401_})
2'b00 : new_n4365_ = 1'b1;
default : new_n4365_ = 1'b0;
endcase
casez ({new_n1111_, new_n1628_})
2'b00 : new_n4366_ = 1'b1;
default : new_n4366_ = 1'b0;
endcase
casez ({new_n80_, new_n1399_, new_n1628_})
3'b01? : new_n4367_ = 1'b1;
3'b??1 : new_n4367_ = 1'b1;
default : new_n4367_ = 1'b0;
endcase
casez ({new_n2646_, new_n3408_})
2'b00 : new_n4368_ = 1'b1;
default : new_n4368_ = 1'b0;
endcase
casez ({new_n2557_, new_n3411_})
2'b00 : new_n4369_ = 1'b1;
default : new_n4369_ = 1'b0;
endcase
casez ({new_n4653_, new_n3414_})
2'b1? : new_n4370_ = 1'b1;
2'b?1 : new_n4370_ = 1'b1;
default : new_n4370_ = 1'b0;
endcase
casez ({new_n1369_, new_n3415_})
2'b00 : new_n4371_ = 1'b1;
default : new_n4371_ = 1'b0;
endcase
casez ({new_n471_, new_n1630_})
2'b00 : new_n4372_ = 1'b1;
default : new_n4372_ = 1'b0;
endcase
casez ({new_n1607_, new_n3420_})
2'b00 : new_n4373_ = 1'b1;
default : new_n4373_ = 1'b0;
endcase
casez ({new_n1863_, new_n3422_})
2'b00 : new_n4374_ = 1'b1;
default : new_n4374_ = 1'b0;
endcase
casez ({new_n1026_, new_n1631_})
2'b00 : new_n4375_ = 1'b1;
default : new_n4375_ = 1'b0;
endcase
casez ({v[2], new_n89_, new_n1035_})
3'b01? : new_n4376_ = 1'b1;
3'b??1 : new_n4376_ = 1'b1;
default : new_n4376_ = 1'b0;
endcase
casez ({new_n2740_, new_n3425_})
2'b00 : new_n4377_ = 1'b1;
default : new_n4377_ = 1'b0;
endcase
casez ({new_n2766_, new_n3426_})
2'b00 : new_n4378_ = 1'b1;
default : new_n4378_ = 1'b0;
endcase
casez ({new_n2556_, new_n3428_})
2'b00 : new_n4379_ = 1'b1;
default : new_n4379_ = 1'b0;
endcase
casez ({new_n659_, new_n1803_, new_n3430_})
3'b01? : new_n4380_ = 1'b1;
3'b??1 : new_n4380_ = 1'b1;
default : new_n4380_ = 1'b0;
endcase
casez ({new_n1143_, new_n3431_})
2'b00 : new_n4381_ = 1'b1;
default : new_n4381_ = 1'b0;
endcase
casez ({new_n158_, new_n398_, new_n178_, new_n309_})
4'b11?? : new_n4382_ = 1'b1;
4'b??11 : new_n4382_ = 1'b1;
default : new_n4382_ = 1'b0;
endcase
casez ({new_n1041_, new_n1633_})
2'b00 : new_n4383_ = 1'b1;
default : new_n4383_ = 1'b0;
endcase
casez ({new_n243_, new_n398_})
2'b00 : new_n4384_ = 1'b1;
default : new_n4384_ = 1'b0;
endcase
casez ({new_n220_, new_n796_, new_n3439_})
3'b11? : new_n4385_ = 1'b1;
3'b??1 : new_n4385_ = 1'b1;
default : new_n4385_ = 1'b0;
endcase
casez ({new_n79_, new_n3440_, new_n1574_})
3'b11? : new_n4386_ = 1'b1;
3'b??1 : new_n4386_ = 1'b1;
default : new_n4386_ = 1'b0;
endcase
casez ({new_n2584_, new_n3443_})
2'b00 : new_n4387_ = 1'b1;
default : new_n4387_ = 1'b0;
endcase
casez ({new_n202_, new_n3445_})
2'b00 : new_n4388_ = 1'b1;
default : new_n4388_ = 1'b0;
endcase
casez ({new_n1633_, new_n3445_})
2'b00 : new_n4389_ = 1'b1;
default : new_n4389_ = 1'b0;
endcase
casez ({new_n435_, new_n1635_})
2'b00 : new_n4390_ = 1'b1;
default : new_n4390_ = 1'b0;
endcase
casez ({new_n2631_, new_n3446_})
2'b00 : new_n4391_ = 1'b1;
default : new_n4391_ = 1'b0;
endcase
casez ({new_n396_, new_n1636_})
2'b00 : new_n4392_ = 1'b1;
default : new_n4392_ = 1'b0;
endcase
casez ({new_n451_, new_n3451_})
2'b00 : new_n4393_ = 1'b1;
default : new_n4393_ = 1'b0;
endcase
casez ({new_n1598_, new_n3453_})
2'b00 : new_n4394_ = 1'b1;
default : new_n4394_ = 1'b0;
endcase
casez ({new_n2673_, new_n3454_})
2'b00 : new_n4395_ = 1'b1;
default : new_n4395_ = 1'b0;
endcase
casez ({new_n323_, new_n1636_})
2'b00 : new_n4396_ = 1'b1;
default : new_n4396_ = 1'b0;
endcase
casez ({new_n1637_, new_n3455_})
2'b00 : new_n4397_ = 1'b1;
default : new_n4397_ = 1'b0;
endcase
casez ({new_n211_, new_n633_, new_n1037_})
3'b11? : new_n4398_ = 1'b1;
3'b??1 : new_n4398_ = 1'b1;
default : new_n4398_ = 1'b0;
endcase
casez ({new_n80_, new_n170_, new_n1638_})
3'b11? : new_n4399_ = 1'b1;
3'b??1 : new_n4399_ = 1'b1;
default : new_n4399_ = 1'b0;
endcase
casez ({new_n788_, new_n3460_})
2'b00 : new_n4400_ = 1'b1;
default : new_n4400_ = 1'b0;
endcase
casez ({new_n1947_, new_n3461_})
2'b00 : new_n4401_ = 1'b1;
default : new_n4401_ = 1'b0;
endcase
casez ({new_n1047_, new_n3465_})
2'b00 : new_n4402_ = 1'b1;
default : new_n4402_ = 1'b0;
endcase
casez ({new_n2675_, new_n3468_})
2'b00 : new_n4403_ = 1'b1;
default : new_n4403_ = 1'b0;
endcase
casez ({new_n1951_, new_n3469_})
2'b00 : new_n4404_ = 1'b1;
default : new_n4404_ = 1'b0;
endcase
casez ({new_n457_, new_n1038_})
2'b00 : new_n4405_ = 1'b1;
default : new_n4405_ = 1'b0;
endcase
casez ({new_n1162_, new_n3472_})
2'b00 : new_n4406_ = 1'b1;
default : new_n4406_ = 1'b0;
endcase
casez ({new_n132_, new_n182_, new_n225_, new_n1039_})
4'b11?? : new_n4407_ = 1'b1;
4'b??11 : new_n4407_ = 1'b1;
default : new_n4407_ = 1'b0;
endcase
casez ({new_n450_, new_n1639_})
2'b00 : new_n4408_ = 1'b1;
default : new_n4408_ = 1'b0;
endcase
casez ({new_n245_, new_n3482_})
2'b00 : new_n4409_ = 1'b1;
default : new_n4409_ = 1'b0;
endcase
casez ({new_n1398_, new_n1640_})
2'b00 : new_n4410_ = 1'b1;
default : new_n4410_ = 1'b0;
endcase
casez ({new_n2575_, new_n3486_})
2'b00 : new_n4411_ = 1'b1;
default : new_n4411_ = 1'b0;
endcase
casez ({new_n1029_, new_n1641_})
2'b00 : new_n4412_ = 1'b1;
default : new_n4412_ = 1'b0;
endcase
casez ({new_n96_, new_n404_, new_n118_, new_n248_})
4'b11?? : new_n4413_ = 1'b1;
4'b??11 : new_n4413_ = 1'b1;
default : new_n4413_ = 1'b0;
endcase
casez ({new_n1160_, new_n1641_})
2'b00 : new_n4414_ = 1'b1;
default : new_n4414_ = 1'b0;
endcase
casez ({new_n795_, new_n1040_})
2'b00 : new_n4415_ = 1'b1;
default : new_n4415_ = 1'b0;
endcase
casez ({new_n536_, new_n1642_})
2'b00 : new_n4416_ = 1'b1;
default : new_n4416_ = 1'b0;
endcase
casez ({new_n421_, new_n3497_})
2'b00 : new_n4417_ = 1'b1;
default : new_n4417_ = 1'b0;
endcase
casez ({new_n104_, new_n1643_, new_n638_})
3'b11? : new_n4418_ = 1'b1;
3'b??1 : new_n4418_ = 1'b1;
default : new_n4418_ = 1'b0;
endcase
casez ({new_n88_, new_n163_, new_n1040_})
3'b01? : new_n4419_ = 1'b1;
3'b??1 : new_n4419_ = 1'b1;
default : new_n4419_ = 1'b0;
endcase
casez ({new_n87_, new_n401_, new_n1644_})
3'b11? : new_n4420_ = 1'b1;
3'b??1 : new_n4420_ = 1'b1;
default : new_n4420_ = 1'b0;
endcase
casez ({new_n311_, new_n405_})
2'b00 : new_n4421_ = 1'b1;
default : new_n4421_ = 1'b0;
endcase
casez ({new_n1558_, new_n3509_})
2'b00 : new_n4422_ = 1'b1;
default : new_n4422_ = 1'b0;
endcase
casez ({new_n336_, new_n3512_})
2'b00 : new_n4423_ = 1'b1;
default : new_n4423_ = 1'b0;
endcase
casez ({new_n345_, new_n1645_})
2'b00 : new_n4424_ = 1'b1;
default : new_n4424_ = 1'b0;
endcase
casez ({new_n737_, new_n3518_})
2'b00 : new_n4425_ = 1'b1;
default : new_n4425_ = 1'b0;
endcase
casez ({new_n1142_, new_n1647_})
2'b00 : new_n4426_ = 1'b1;
default : new_n4426_ = 1'b0;
endcase
casez ({new_n1646_, new_n3528_})
2'b00 : new_n4427_ = 1'b1;
default : new_n4427_ = 1'b0;
endcase
casez ({new_n2754_, new_n3529_})
2'b00 : new_n4428_ = 1'b1;
default : new_n4428_ = 1'b0;
endcase
casez ({new_n153_, new_n393_, new_n3536_})
3'b10? : new_n4429_ = 1'b1;
3'b??1 : new_n4429_ = 1'b1;
default : new_n4429_ = 1'b0;
endcase
casez ({new_n1578_, new_n1648_})
2'b00 : new_n4430_ = 1'b1;
default : new_n4430_ = 1'b0;
endcase
casez ({new_n2632_, new_n3538_})
2'b00 : new_n4431_ = 1'b1;
default : new_n4431_ = 1'b0;
endcase
casez ({new_n1028_, new_n1649_})
2'b00 : new_n4432_ = 1'b1;
default : new_n4432_ = 1'b0;
endcase
casez ({new_n258_, new_n358_, new_n1043_})
3'b11? : new_n4433_ = 1'b1;
3'b??1 : new_n4433_ = 1'b1;
default : new_n4433_ = 1'b0;
endcase
casez ({new_n4622_, new_n107_, new_n124_})
3'b1?? : new_n4434_ = 1'b1;
3'b?01 : new_n4434_ = 1'b1;
default : new_n4434_ = 1'b0;
endcase
casez ({new_n1931_, new_n3542_})
2'b00 : new_n4435_ = 1'b1;
default : new_n4435_ = 1'b0;
endcase
casez ({new_n2687_, new_n3546_})
2'b00 : new_n4436_ = 1'b1;
default : new_n4436_ = 1'b0;
endcase
casez ({new_n740_, new_n3546_})
2'b00 : new_n4437_ = 1'b1;
default : new_n4437_ = 1'b0;
endcase
casez ({new_n2637_, new_n3550_})
2'b00 : new_n4438_ = 1'b1;
default : new_n4438_ = 1'b0;
endcase
casez ({new_n93_, new_n3552_, new_n619_, new_n1867_})
4'b01?? : new_n4439_ = 1'b1;
4'b??11 : new_n4439_ = 1'b1;
default : new_n4439_ = 1'b0;
endcase
casez ({new_n92_, new_n3553_, new_n1842_})
3'b11? : new_n4440_ = 1'b1;
3'b??1 : new_n4440_ = 1'b1;
default : new_n4440_ = 1'b0;
endcase
casez ({new_n494_, new_n3558_})
2'b00 : new_n4441_ = 1'b1;
default : new_n4441_ = 1'b0;
endcase
casez ({new_n1651_, new_n3564_})
2'b00 : new_n4442_ = 1'b1;
default : new_n4442_ = 1'b0;
endcase
casez ({new_n455_, new_n3565_})
2'b00 : new_n4443_ = 1'b1;
default : new_n4443_ = 1'b0;
endcase
casez ({new_n1402_, new_n3566_})
2'b00 : new_n4444_ = 1'b1;
default : new_n4444_ = 1'b0;
endcase
casez ({new_n245_, new_n3567_})
2'b00 : new_n4445_ = 1'b1;
default : new_n4445_ = 1'b0;
endcase
casez ({new_n83_, new_n152_, new_n1046_})
3'b11? : new_n4446_ = 1'b1;
3'b??1 : new_n4446_ = 1'b1;
default : new_n4446_ = 1'b0;
endcase
casez ({new_n671_, new_n3571_})
2'b00 : new_n4447_ = 1'b1;
default : new_n4447_ = 1'b0;
endcase
casez ({new_n391_, new_n3572_})
2'b00 : new_n4448_ = 1'b1;
default : new_n4448_ = 1'b0;
endcase
casez ({new_n1126_, new_n3578_})
2'b00 : new_n4449_ = 1'b1;
default : new_n4449_ = 1'b0;
endcase
casez ({new_n1370_, new_n3582_})
2'b00 : new_n4450_ = 1'b1;
default : new_n4450_ = 1'b0;
endcase
casez ({new_n350_, new_n3586_})
2'b00 : new_n4451_ = 1'b1;
default : new_n4451_ = 1'b0;
endcase
casez ({v[0], new_n1045_, new_n333_, new_n396_})
4'b01?? : new_n4452_ = 1'b1;
4'b??01 : new_n4452_ = 1'b1;
default : new_n4452_ = 1'b0;
endcase
casez ({new_n185_, new_n3588_})
2'b00 : new_n4453_ = 1'b1;
default : new_n4453_ = 1'b0;
endcase
casez ({new_n100_, new_n3596_, new_n1146_})
3'b01? : new_n4454_ = 1'b1;
3'b??1 : new_n4454_ = 1'b1;
default : new_n4454_ = 1'b0;
endcase
casez ({new_n2732_, new_n3597_})
2'b00 : new_n4455_ = 1'b1;
default : new_n4455_ = 1'b0;
endcase
casez ({new_n525_, new_n3598_})
2'b00 : new_n4456_ = 1'b1;
default : new_n4456_ = 1'b0;
endcase
casez ({new_n220_, new_n398_, new_n710_})
3'b11? : new_n4457_ = 1'b1;
3'b??1 : new_n4457_ = 1'b1;
default : new_n4457_ = 1'b0;
endcase
casez ({new_n1827_, new_n3604_})
2'b00 : new_n4458_ = 1'b1;
default : new_n4458_ = 1'b0;
endcase
casez ({new_n179_, new_n209_, new_n710_})
3'b11? : new_n4459_ = 1'b1;
3'b??1 : new_n4459_ = 1'b1;
default : new_n4459_ = 1'b0;
endcase
casez ({new_n247_, new_n302_, new_n711_})
3'b10? : new_n4460_ = 1'b1;
3'b??1 : new_n4460_ = 1'b1;
default : new_n4460_ = 1'b0;
endcase
casez ({new_n154_, new_n712_})
2'b00 : new_n4461_ = 1'b1;
default : new_n4461_ = 1'b0;
endcase
casez ({new_n86_, new_n712_, new_n104_, new_n541_})
4'b11?? : new_n4462_ = 1'b1;
4'b??11 : new_n4462_ = 1'b1;
default : new_n4462_ = 1'b0;
endcase
casez ({new_n584_, new_n713_})
2'b00 : new_n4463_ = 1'b1;
default : new_n4463_ = 1'b0;
endcase
casez ({new_n334_, new_n713_})
2'b00 : new_n4464_ = 1'b1;
default : new_n4464_ = 1'b0;
endcase
casez ({new_n80_, new_n176_, new_n714_})
3'b11? : new_n4465_ = 1'b1;
3'b??1 : new_n4465_ = 1'b1;
default : new_n4465_ = 1'b0;
endcase
casez ({new_n538_, new_n716_})
2'b00 : new_n4466_ = 1'b1;
default : new_n4466_ = 1'b0;
endcase
casez ({new_n265_, new_n716_})
2'b00 : new_n4467_ = 1'b1;
default : new_n4467_ = 1'b0;
endcase
casez ({new_n185_, new_n421_})
2'b00 : new_n4468_ = 1'b1;
default : new_n4468_ = 1'b0;
endcase
casez ({new_n250_, new_n422_, new_n299_, new_n398_})
4'b11?? : new_n4469_ = 1'b1;
4'b??11 : new_n4469_ = 1'b1;
default : new_n4469_ = 1'b0;
endcase
casez ({new_n94_, new_n115_, new_n260_, new_n422_})
4'b11?? : new_n4470_ = 1'b1;
4'b??11 : new_n4470_ = 1'b1;
default : new_n4470_ = 1'b0;
endcase
casez ({new_n671_, new_n718_})
2'b00 : new_n4471_ = 1'b1;
default : new_n4471_ = 1'b0;
endcase
casez ({new_n451_, new_n718_})
2'b00 : new_n4472_ = 1'b1;
default : new_n4472_ = 1'b0;
endcase
casez ({new_n243_, new_n719_})
2'b00 : new_n4473_ = 1'b1;
default : new_n4473_ = 1'b0;
endcase
casez ({new_n81_, new_n429_, new_n316_, new_n352_})
4'b11?? : new_n4474_ = 1'b1;
4'b??11 : new_n4474_ = 1'b1;
default : new_n4474_ = 1'b0;
endcase
casez ({new_n282_, new_n441_})
2'b00 : new_n4475_ = 1'b1;
default : new_n4475_ = 1'b0;
endcase
casez ({new_n85_, new_n257_, new_n441_})
3'b11? : new_n4476_ = 1'b1;
3'b??1 : new_n4476_ = 1'b1;
default : new_n4476_ = 1'b0;
endcase
casez ({new_n236_, new_n1098_})
2'b00 : new_n4477_ = 1'b1;
default : new_n4477_ = 1'b0;
endcase
casez ({new_n711_, new_n735_})
2'b00 : new_n4478_ = 1'b1;
default : new_n4478_ = 1'b0;
endcase
casez ({new_n864_, new_n1099_})
2'b00 : new_n4479_ = 1'b1;
default : new_n4479_ = 1'b0;
endcase
casez ({x[2], new_n1103_, new_n95_, new_n183_})
4'b11?? : new_n4480_ = 1'b1;
4'b??11 : new_n4480_ = 1'b1;
default : new_n4480_ = 1'b0;
endcase
casez ({new_n960_, new_n1799_})
2'b00 : new_n4481_ = 1'b1;
default : new_n4481_ = 1'b0;
endcase
casez ({new_n387_, new_n1800_})
2'b00 : new_n4482_ = 1'b1;
default : new_n4482_ = 1'b0;
endcase
casez ({new_n1344_, new_n1800_})
2'b00 : new_n4483_ = 1'b1;
default : new_n4483_ = 1'b0;
endcase
casez ({new_n1583_, new_n1800_})
2'b00 : new_n4484_ = 1'b1;
default : new_n4484_ = 1'b0;
endcase
casez ({new_n527_, new_n737_})
2'b00 : new_n4485_ = 1'b1;
default : new_n4485_ = 1'b0;
endcase
casez ({new_n104_, new_n728_, new_n1107_})
3'b11? : new_n4486_ = 1'b1;
3'b??1 : new_n4486_ = 1'b1;
default : new_n4486_ = 1'b0;
endcase
casez ({new_n310_, new_n1107_})
2'b00 : new_n4487_ = 1'b1;
default : new_n4487_ = 1'b0;
endcase
casez ({new_n710_, new_n738_})
2'b00 : new_n4488_ = 1'b1;
default : new_n4488_ = 1'b0;
endcase
casez ({new_n186_, new_n207_, new_n738_})
3'b11? : new_n4489_ = 1'b1;
3'b??1 : new_n4489_ = 1'b1;
default : new_n4489_ = 1'b0;
endcase
casez ({new_n710_, new_n1109_})
2'b00 : new_n4490_ = 1'b1;
default : new_n4490_ = 1'b0;
endcase
casez ({new_n194_, new_n420_, new_n1109_})
3'b11? : new_n4491_ = 1'b1;
3'b??1 : new_n4491_ = 1'b1;
default : new_n4491_ = 1'b0;
endcase
casez ({new_n310_, new_n455_})
2'b00 : new_n4492_ = 1'b1;
default : new_n4492_ = 1'b0;
endcase
casez ({new_n1042_, new_n1110_})
2'b00 : new_n4493_ = 1'b1;
default : new_n4493_ = 1'b0;
endcase
casez ({new_n144_, new_n219_, new_n1111_})
3'b11? : new_n4494_ = 1'b1;
3'b??1 : new_n4494_ = 1'b1;
default : new_n4494_ = 1'b0;
endcase
casez ({x[1], new_n259_, new_n1111_})
3'b01? : new_n4495_ = 1'b1;
3'b??1 : new_n4495_ = 1'b1;
default : new_n4495_ = 1'b0;
endcase
casez ({new_n4666_, new_n113_, new_n115_})
3'b1?? : new_n4496_ = 1'b1;
3'b?11 : new_n4496_ = 1'b1;
default : new_n4496_ = 1'b0;
endcase
casez ({new_n112_, new_n183_, new_n1822_})
3'b11? : new_n4497_ = 1'b1;
3'b??1 : new_n4497_ = 1'b1;
default : new_n4497_ = 1'b0;
endcase
casez ({new_n159_, new_n252_, new_n1822_})
3'b10? : new_n4498_ = 1'b1;
3'b??1 : new_n4498_ = 1'b1;
default : new_n4498_ = 1'b0;
endcase
casez ({new_n441_, new_n1823_})
2'b00 : new_n4499_ = 1'b1;
default : new_n4499_ = 1'b0;
endcase
casez ({new_n1589_, new_n1824_})
2'b00 : new_n4500_ = 1'b1;
default : new_n4500_ = 1'b0;
endcase
casez ({new_n581_, new_n1824_})
2'b00 : new_n4501_ = 1'b1;
default : new_n4501_ = 1'b0;
endcase
casez ({new_n1590_, new_n1824_})
2'b00 : new_n4502_ = 1'b1;
default : new_n4502_ = 1'b0;
endcase
casez ({new_n861_, new_n1825_})
2'b00 : new_n4503_ = 1'b1;
default : new_n4503_ = 1'b0;
endcase
casez ({new_n940_, new_n1113_})
2'b00 : new_n4504_ = 1'b1;
default : new_n4504_ = 1'b0;
endcase
casez ({y[2], new_n454_, new_n83_, new_n1113_})
4'b01?? : new_n4505_ = 1'b1;
4'b??01 : new_n4505_ = 1'b1;
default : new_n4505_ = 1'b0;
endcase
casez ({new_n95_, new_n147_, new_n460_})
3'b01? : new_n4506_ = 1'b1;
3'b??1 : new_n4506_ = 1'b1;
default : new_n4506_ = 1'b0;
endcase
casez ({new_n171_, new_n460_})
2'b00 : new_n4507_ = 1'b1;
default : new_n4507_ = 1'b0;
endcase
casez ({new_n200_, new_n338_, new_n1115_})
3'b11? : new_n4508_ = 1'b1;
3'b??1 : new_n4508_ = 1'b1;
default : new_n4508_ = 1'b0;
endcase
casez ({new_n139_, new_n413_, new_n1831_})
3'b10? : new_n4509_ = 1'b1;
3'b??1 : new_n4509_ = 1'b1;
default : new_n4509_ = 1'b0;
endcase
casez ({new_n386_, new_n460_})
2'b00 : new_n4510_ = 1'b1;
default : new_n4510_ = 1'b0;
endcase
casez ({new_n166_, new_n358_, new_n1833_})
3'b11? : new_n4511_ = 1'b1;
3'b??1 : new_n4511_ = 1'b1;
default : new_n4511_ = 1'b0;
endcase
casez ({new_n1364_, new_n1833_})
2'b00 : new_n4512_ = 1'b1;
default : new_n4512_ = 1'b0;
endcase
casez ({new_n718_, new_n1114_})
2'b00 : new_n4513_ = 1'b1;
default : new_n4513_ = 1'b0;
endcase
casez ({new_n208_, new_n469_, new_n1117_})
3'b11? : new_n4514_ = 1'b1;
3'b??1 : new_n4514_ = 1'b1;
default : new_n4514_ = 1'b0;
endcase
casez ({u[2], new_n681_, new_n1836_})
3'b11? : new_n4515_ = 1'b1;
3'b??1 : new_n4515_ = 1'b1;
default : new_n4515_ = 1'b0;
endcase
casez ({new_n1027_, new_n1118_})
2'b00 : new_n4516_ = 1'b1;
default : new_n4516_ = 1'b0;
endcase
casez ({new_n4634_, new_n1840_})
2'b1? : new_n4517_ = 1'b1;
2'b?1 : new_n4517_ = 1'b1;
default : new_n4517_ = 1'b0;
endcase
casez ({new_n196_, new_n541_, new_n1840_})
3'b11? : new_n4518_ = 1'b1;
3'b??1 : new_n4518_ = 1'b1;
default : new_n4518_ = 1'b0;
endcase
casez ({new_n1639_, new_n1841_})
2'b00 : new_n4519_ = 1'b1;
default : new_n4519_ = 1'b0;
endcase
casez ({new_n319_, new_n451_, new_n1120_})
3'b01? : new_n4520_ = 1'b1;
3'b??1 : new_n4520_ = 1'b1;
default : new_n4520_ = 1'b0;
endcase
casez ({new_n1569_, new_n1845_})
2'b00 : new_n4521_ = 1'b1;
default : new_n4521_ = 1'b0;
endcase
casez ({new_n1167_, new_n1846_})
2'b00 : new_n4522_ = 1'b1;
default : new_n4522_ = 1'b0;
endcase
casez ({new_n89_, new_n383_, new_n1847_})
3'b11? : new_n4523_ = 1'b1;
3'b??1 : new_n4523_ = 1'b1;
default : new_n4523_ = 1'b0;
endcase
casez ({new_n4637_, new_n367_})
2'b1? : new_n4524_ = 1'b1;
2'b?1 : new_n4524_ = 1'b1;
default : new_n4524_ = 1'b0;
endcase
casez ({new_n82_, new_n192_, new_n1849_})
3'b11? : new_n4525_ = 1'b1;
3'b??1 : new_n4525_ = 1'b1;
default : new_n4525_ = 1'b0;
endcase
casez ({new_n1026_, new_n1124_})
2'b00 : new_n4526_ = 1'b1;
default : new_n4526_ = 1'b0;
endcase
casez ({new_n150_, new_n318_, new_n1853_})
3'b11? : new_n4527_ = 1'b1;
3'b??1 : new_n4527_ = 1'b1;
default : new_n4527_ = 1'b0;
endcase
casez ({new_n1122_, new_n1853_})
2'b00 : new_n4528_ = 1'b1;
default : new_n4528_ = 1'b0;
endcase
casez ({new_n1594_, new_n1854_})
2'b00 : new_n4529_ = 1'b1;
default : new_n4529_ = 1'b0;
endcase
casez ({new_n178_, new_n1125_})
2'b00 : new_n4530_ = 1'b1;
default : new_n4530_ = 1'b0;
endcase
casez ({new_n1144_, new_n1855_})
2'b00 : new_n4531_ = 1'b1;
default : new_n4531_ = 1'b0;
endcase
casez ({u[2], new_n187_, new_n1125_})
3'b11? : new_n4532_ = 1'b1;
3'b??1 : new_n4532_ = 1'b1;
default : new_n4532_ = 1'b0;
endcase
casez ({new_n677_, new_n1856_})
2'b00 : new_n4533_ = 1'b1;
default : new_n4533_ = 1'b0;
endcase
casez ({new_n347_, new_n1125_})
2'b00 : new_n4534_ = 1'b1;
default : new_n4534_ = 1'b0;
endcase
casez ({new_n334_, new_n1126_})
2'b00 : new_n4535_ = 1'b1;
default : new_n4535_ = 1'b0;
endcase
casez ({new_n1014_, new_n1858_})
2'b00 : new_n4536_ = 1'b1;
default : new_n4536_ = 1'b0;
endcase
casez ({new_n1007_, new_n1860_})
2'b00 : new_n4537_ = 1'b1;
default : new_n4537_ = 1'b0;
endcase
casez ({new_n471_, new_n1863_})
2'b00 : new_n4538_ = 1'b1;
default : new_n4538_ = 1'b0;
endcase
casez ({new_n767_, new_n1863_})
2'b00 : new_n4539_ = 1'b1;
default : new_n4539_ = 1'b0;
endcase
casez ({new_n1030_, new_n1864_})
2'b00 : new_n4540_ = 1'b1;
default : new_n4540_ = 1'b0;
endcase
casez ({new_n1558_, new_n1865_})
2'b00 : new_n4541_ = 1'b1;
default : new_n4541_ = 1'b0;
endcase
casez ({new_n1266_, new_n1866_})
2'b00 : new_n4542_ = 1'b1;
default : new_n4542_ = 1'b0;
endcase
casez ({new_n1147_, new_n1868_})
2'b00 : new_n4543_ = 1'b1;
default : new_n4543_ = 1'b0;
endcase
casez ({new_n1351_, new_n1870_})
2'b00 : new_n4544_ = 1'b1;
default : new_n4544_ = 1'b0;
endcase
casez ({new_n176_, new_n275_, new_n1870_})
3'b11? : new_n4545_ = 1'b1;
3'b??1 : new_n4545_ = 1'b1;
default : new_n4545_ = 1'b0;
endcase
casez ({new_n859_, new_n1131_})
2'b00 : new_n4546_ = 1'b1;
default : new_n4546_ = 1'b0;
endcase
casez ({new_n740_, new_n1131_})
2'b00 : new_n4547_ = 1'b1;
default : new_n4547_ = 1'b0;
endcase
casez ({new_n1572_, new_n1875_})
2'b00 : new_n4548_ = 1'b1;
default : new_n4548_ = 1'b0;
endcase
casez ({new_n1144_, new_n1875_})
2'b00 : new_n4549_ = 1'b1;
default : new_n4549_ = 1'b0;
endcase
casez ({new_n752_, new_n1133_})
2'b00 : new_n4550_ = 1'b1;
default : new_n4550_ = 1'b0;
endcase
casez ({new_n503_, new_n1134_})
2'b00 : new_n4551_ = 1'b1;
default : new_n4551_ = 1'b0;
endcase
casez ({new_n383_, new_n438_, new_n1878_})
3'b11? : new_n4552_ = 1'b1;
3'b??1 : new_n4552_ = 1'b1;
default : new_n4552_ = 1'b0;
endcase
casez ({new_n1826_, new_n1879_})
2'b00 : new_n4553_ = 1'b1;
default : new_n4553_ = 1'b0;
endcase
casez ({v[1], new_n239_, new_n1880_})
3'b01? : new_n4554_ = 1'b1;
3'b??1 : new_n4554_ = 1'b1;
default : new_n4554_ = 1'b0;
endcase
casez ({u[2], new_n301_, new_n1134_})
3'b01? : new_n4555_ = 1'b1;
3'b??1 : new_n4555_ = 1'b1;
default : new_n4555_ = 1'b0;
endcase
casez ({new_n173_, new_n1881_})
2'b00 : new_n4556_ = 1'b1;
default : new_n4556_ = 1'b0;
endcase
casez ({new_n142_, new_n1882_, new_n378_, new_n398_})
4'b11?? : new_n4557_ = 1'b1;
4'b??11 : new_n4557_ = 1'b1;
default : new_n4557_ = 1'b0;
endcase
casez ({new_n85_, new_n1882_, new_n106_, new_n201_})
4'b11?? : new_n4558_ = 1'b1;
4'b??11 : new_n4558_ = 1'b1;
default : new_n4558_ = 1'b0;
endcase
casez ({new_n4591_, new_n1136_})
2'b1? : new_n4559_ = 1'b1;
2'b?1 : new_n4559_ = 1'b1;
default : new_n4559_ = 1'b0;
endcase
casez ({x[0], new_n1884_, new_n1364_})
3'b01? : new_n4560_ = 1'b1;
3'b??1 : new_n4560_ = 1'b1;
default : new_n4560_ = 1'b0;
endcase
casez ({new_n1837_, new_n1886_})
2'b00 : new_n4561_ = 1'b1;
default : new_n4561_ = 1'b0;
endcase
casez ({new_n158_, new_n207_, new_n1139_})
3'b11? : new_n4562_ = 1'b1;
3'b??1 : new_n4562_ = 1'b1;
default : new_n4562_ = 1'b0;
endcase
casez ({new_n182_, new_n491_, new_n1890_})
3'b10? : new_n4563_ = 1'b1;
3'b??1 : new_n4563_ = 1'b1;
default : new_n4563_ = 1'b0;
endcase
casez ({new_n1138_, new_n1139_})
2'b00 : new_n4564_ = 1'b1;
default : new_n4564_ = 1'b0;
endcase
casez ({new_n869_, new_n1893_})
2'b00 : new_n4565_ = 1'b1;
default : new_n4565_ = 1'b0;
endcase
casez ({new_n273_, new_n302_, new_n1896_})
3'b10? : new_n4566_ = 1'b1;
3'b??1 : new_n4566_ = 1'b1;
default : new_n4566_ = 1'b0;
endcase
casez ({new_n1618_, new_n1896_})
2'b00 : new_n4567_ = 1'b1;
default : new_n4567_ = 1'b0;
endcase
casez ({new_n1106_, new_n1897_})
2'b00 : new_n4568_ = 1'b1;
default : new_n4568_ = 1'b0;
endcase
casez ({new_n4634_, new_n1142_})
2'b1? : new_n4569_ = 1'b1;
2'b?1 : new_n4569_ = 1'b1;
default : new_n4569_ = 1'b0;
endcase
casez ({new_n1348_, new_n1900_})
2'b00 : new_n4570_ = 1'b1;
default : new_n4570_ = 1'b0;
endcase
casez ({y[2], new_n503_, new_n153_, new_n200_})
4'b11?? : new_n4571_ = 1'b1;
4'b??11 : new_n4571_ = 1'b1;
default : new_n4571_ = 1'b0;
endcase
casez ({new_n286_, new_n504_})
2'b00 : new_n4572_ = 1'b1;
default : new_n4572_ = 1'b0;
endcase
casez ({new_n185_, new_n286_})
2'b00 : new_n4573_ = 1'b1;
default : new_n4573_ = 1'b0;
endcase
casez ({new_n121_, new_n333_})
2'b01 : new_n4574_ = 1'b1;
default : new_n4574_ = 1'b0;
endcase
casez ({new_n126_, new_n336_})
2'b00 : new_n4575_ = 1'b1;
default : new_n4575_ = 1'b0;
endcase
casez ({new_n94_, new_n101_, new_n372_})
3'b11? : new_n4576_ = 1'b1;
3'b??1 : new_n4576_ = 1'b1;
default : new_n4576_ = 1'b0;
endcase
casez ({new_n115_, new_n430_})
2'b00 : new_n4577_ = 1'b1;
default : new_n4577_ = 1'b0;
endcase
casez ({new_n88_, new_n127_, new_n89_, new_n106_})
4'b11?? : new_n4578_ = 1'b1;
4'b??11 : new_n4578_ = 1'b1;
default : new_n4578_ = 1'b0;
endcase
casez ({new_n284_, new_n465_})
2'b01 : new_n4579_ = 1'b1;
default : new_n4579_ = 1'b0;
endcase
casez ({new_n77_, new_n483_})
2'b01 : new_n4580_ = 1'b1;
default : new_n4580_ = 1'b0;
endcase
casez ({new_n511_, new_n1151_})
2'b01 : new_n4581_ = 1'b1;
default : new_n4581_ = 1'b0;
endcase
casez ({new_n201_, new_n778_})
2'b11 : new_n4582_ = 1'b1;
default : new_n4582_ = 1'b0;
endcase
casez ({u[0], new_n781_})
2'b01 : new_n4583_ = 1'b1;
default : new_n4583_ = 1'b0;
endcase
casez ({new_n158_, new_n784_})
2'b11 : new_n4584_ = 1'b1;
default : new_n4584_ = 1'b0;
endcase
casez ({x[0], new_n781_})
2'b11 : new_n4585_ = 1'b1;
default : new_n4585_ = 1'b0;
endcase
casez ({new_n632_, new_n1173_})
2'b11 : new_n4586_ = 1'b1;
default : new_n4586_ = 1'b0;
endcase
casez ({new_n96_, new_n790_})
2'b11 : new_n4587_ = 1'b1;
default : new_n4587_ = 1'b0;
endcase
casez ({y[0], new_n526_})
2'b11 : new_n4588_ = 1'b1;
default : new_n4588_ = 1'b0;
endcase
casez ({new_n85_, new_n537_})
2'b11 : new_n4589_ = 1'b1;
default : new_n4589_ = 1'b0;
endcase
casez ({new_n238_, new_n541_})
2'b11 : new_n4590_ = 1'b1;
default : new_n4590_ = 1'b0;
endcase
casez ({u[0], new_n543_})
2'b11 : new_n4591_ = 1'b1;
default : new_n4591_ = 1'b0;
endcase
casez ({new_n148_, new_n1296_})
2'b10 : new_n4592_ = 1'b1;
default : new_n4592_ = 1'b0;
endcase
casez ({new_n89_, new_n294_})
2'b01 : new_n4593_ = 1'b1;
default : new_n4593_ = 1'b0;
endcase
casez ({new_n476_, new_n580_})
2'b11 : new_n4594_ = 1'b1;
default : new_n4594_ = 1'b0;
endcase
casez ({new_n261_, new_n1350_})
2'b11 : new_n4595_ = 1'b1;
default : new_n4595_ = 1'b0;
endcase
casez ({new_n228_, new_n1350_})
2'b11 : new_n4596_ = 1'b1;
default : new_n4596_ = 1'b0;
endcase
casez ({x[0], new_n583_})
2'b11 : new_n4597_ = 1'b1;
default : new_n4597_ = 1'b0;
endcase
casez ({u[0], new_n581_})
2'b11 : new_n4598_ = 1'b1;
default : new_n4598_ = 1'b0;
endcase
casez ({new_n97_, new_n320_})
2'b10 : new_n4599_ = 1'b1;
default : new_n4599_ = 1'b0;
endcase
casez ({new_n360_, new_n2589_})
2'b11 : new_n4600_ = 1'b1;
default : new_n4600_ = 1'b0;
endcase
casez ({new_n214_, new_n935_})
2'b10 : new_n4601_ = 1'b1;
default : new_n4601_ = 1'b0;
endcase
casez ({u[0], new_n2639_})
2'b11 : new_n4602_ = 1'b1;
default : new_n4602_ = 1'b0;
endcase
casez ({new_n85_, new_n632_})
2'b01 : new_n4603_ = 1'b1;
default : new_n4603_ = 1'b0;
endcase
casez ({x[0], new_n950_})
2'b01 : new_n4604_ = 1'b1;
default : new_n4604_ = 1'b0;
endcase
casez ({y[1], new_n961_})
2'b11 : new_n4605_ = 1'b1;
default : new_n4605_ = 1'b0;
endcase
casez ({new_n114_, new_n352_})
2'b11 : new_n4606_ = 1'b1;
default : new_n4606_ = 1'b0;
endcase
casez ({new_n157_, new_n363_})
2'b11 : new_n4607_ = 1'b1;
default : new_n4607_ = 1'b0;
endcase
casez ({new_n472_, new_n2971_})
2'b11 : new_n4608_ = 1'b1;
default : new_n4608_ = 1'b0;
endcase
casez ({new_n119_, new_n372_})
2'b11 : new_n4609_ = 1'b1;
default : new_n4609_ = 1'b0;
endcase
casez ({v[0], new_n102_})
2'b11 : new_n4610_ = 1'b1;
default : new_n4610_ = 1'b0;
endcase
casez ({new_n91_, new_n1005_})
2'b11 : new_n4611_ = 1'b1;
default : new_n4611_ = 1'b0;
endcase
casez ({u[0], new_n382_})
2'b11 : new_n4612_ = 1'b1;
default : new_n4612_ = 1'b0;
endcase
casez ({new_n100_, new_n680_})
2'b11 : new_n4613_ = 1'b1;
default : new_n4613_ = 1'b0;
endcase
casez ({new_n229_, new_n388_})
2'b11 : new_n4614_ = 1'b1;
default : new_n4614_ = 1'b0;
endcase
casez ({new_n86_, new_n387_})
2'b01 : new_n4615_ = 1'b1;
default : new_n4615_ = 1'b0;
endcase
casez ({v[0], new_n1613_})
2'b01 : new_n4616_ = 1'b1;
default : new_n4616_ = 1'b0;
endcase
casez ({new_n88_, new_n390_})
2'b11 : new_n4617_ = 1'b1;
default : new_n4617_ = 1'b0;
endcase
casez ({new_n476_, new_n3360_})
2'b11 : new_n4618_ = 1'b1;
default : new_n4618_ = 1'b0;
endcase
casez ({new_n77_, new_n395_})
2'b01 : new_n4619_ = 1'b1;
default : new_n4619_ = 1'b0;
endcase
casez ({new_n243_, new_n395_})
2'b11 : new_n4620_ = 1'b1;
default : new_n4620_ = 1'b0;
endcase
casez ({new_n80_, new_n1650_})
2'b01 : new_n4621_ = 1'b1;
default : new_n4621_ = 1'b0;
endcase
casez ({u[2], new_n408_})
2'b01 : new_n4622_ = 1'b1;
default : new_n4622_ = 1'b0;
endcase
casez ({new_n183_, new_n1044_})
2'b11 : new_n4623_ = 1'b1;
default : new_n4623_ = 1'b0;
endcase
casez ({new_n317_, new_n420_})
2'b11 : new_n4624_ = 1'b1;
default : new_n4624_ = 1'b0;
endcase
casez ({new_n235_, new_n430_})
2'b11 : new_n4625_ = 1'b1;
default : new_n4625_ = 1'b0;
endcase
casez ({new_n77_, new_n449_})
2'b01 : new_n4626_ = 1'b1;
default : new_n4626_ = 1'b0;
endcase
casez ({v[2], new_n449_})
2'b11 : new_n4627_ = 1'b1;
default : new_n4627_ = 1'b0;
endcase
casez ({new_n199_, new_n1104_})
2'b11 : new_n4628_ = 1'b1;
default : new_n4628_ = 1'b0;
endcase
casez ({new_n89_, new_n455_})
2'b11 : new_n4629_ = 1'b1;
default : new_n4629_ = 1'b0;
endcase
casez ({new_n88_, new_n455_})
2'b01 : new_n4630_ = 1'b1;
default : new_n4630_ = 1'b0;
endcase
casez ({new_n79_, new_n456_})
2'b01 : new_n4631_ = 1'b1;
default : new_n4631_ = 1'b0;
endcase
casez ({new_n105_, new_n741_})
2'b11 : new_n4632_ = 1'b1;
default : new_n4632_ = 1'b0;
endcase
casez ({x[0], new_n459_})
2'b11 : new_n4633_ = 1'b1;
default : new_n4633_ = 1'b0;
endcase
casez ({u[0], new_n459_})
2'b11 : new_n4634_ = 1'b1;
default : new_n4634_ = 1'b0;
endcase
casez ({new_n154_, new_n1843_})
2'b11 : new_n4635_ = 1'b1;
default : new_n4635_ = 1'b0;
endcase
casez ({new_n542_, new_n750_})
2'b11 : new_n4636_ = 1'b1;
default : new_n4636_ = 1'b0;
endcase
casez ({x[0], new_n749_})
2'b11 : new_n4637_ = 1'b1;
default : new_n4637_ = 1'b0;
endcase
casez ({new_n237_, new_n1852_})
2'b11 : new_n4638_ = 1'b1;
default : new_n4638_ = 1'b0;
endcase
casez ({new_n319_, new_n1131_})
2'b01 : new_n4639_ = 1'b1;
default : new_n4639_ = 1'b0;
endcase
casez ({new_n1025_, new_n1937_})
2'b11 : new_n4640_ = 1'b1;
default : new_n4640_ = 1'b0;
endcase
casez ({new_n93_, new_n259_})
2'b11 : new_n4641_ = 1'b1;
default : new_n4641_ = 1'b0;
endcase
casez ({u[0], new_n517_})
2'b11 : new_n4642_ = 1'b1;
default : new_n4642_ = 1'b0;
endcase
casez ({new_n138_, new_n535_})
2'b11 : new_n4643_ = 1'b1;
default : new_n4643_ = 1'b0;
endcase
casez ({y[2], new_n286_})
2'b11 : new_n4644_ = 1'b1;
default : new_n4644_ = 1'b0;
endcase
casez ({new_n133_, new_n558_})
2'b11 : new_n4645_ = 1'b1;
default : new_n4645_ = 1'b0;
endcase
casez ({new_n223_, new_n619_})
2'b11 : new_n4646_ = 1'b1;
default : new_n4646_ = 1'b0;
endcase
casez ({new_n148_, new_n631_})
2'b11 : new_n4647_ = 1'b1;
default : new_n4647_ = 1'b0;
endcase
casez ({new_n97_, new_n352_})
2'b11 : new_n4648_ = 1'b1;
default : new_n4648_ = 1'b0;
endcase
casez ({new_n119_, new_n202_})
2'b11 : new_n4649_ = 1'b1;
default : new_n4649_ = 1'b0;
endcase
casez ({new_n98_, new_n360_})
2'b11 : new_n4650_ = 1'b1;
default : new_n4650_ = 1'b0;
endcase
casez ({v[1], new_n362_})
2'b01 : new_n4651_ = 1'b1;
default : new_n4651_ = 1'b0;
endcase
casez ({x[0], new_n669_})
2'b11 : new_n4652_ = 1'b1;
default : new_n4652_ = 1'b0;
endcase
casez ({new_n101_, new_n671_})
2'b11 : new_n4653_ = 1'b1;
default : new_n4653_ = 1'b0;
endcase
casez ({new_n84_, new_n380_})
2'b10 : new_n4654_ = 1'b1;
default : new_n4654_ = 1'b0;
endcase
casez ({new_n83_, new_n381_})
2'b11 : new_n4655_ = 1'b1;
default : new_n4655_ = 1'b0;
endcase
casez ({new_n96_, new_n382_})
2'b11 : new_n4656_ = 1'b1;
default : new_n4656_ = 1'b0;
endcase
casez ({x[0], new_n383_})
2'b11 : new_n4657_ = 1'b1;
default : new_n4657_ = 1'b0;
endcase
casez ({new_n85_, new_n389_})
2'b11 : new_n4658_ = 1'b1;
default : new_n4658_ = 1'b0;
endcase
casez ({y[2], new_n393_})
2'b10 : new_n4659_ = 1'b1;
default : new_n4659_ = 1'b0;
endcase
casez ({new_n159_, new_n1032_})
2'b11 : new_n4660_ = 1'b1;
default : new_n4660_ = 1'b0;
endcase
casez ({new_n279_, new_n419_})
2'b11 : new_n4661_ = 1'b1;
default : new_n4661_ = 1'b0;
endcase
casez ({y[2], new_n424_})
2'b11 : new_n4662_ = 1'b1;
default : new_n4662_ = 1'b0;
endcase
casez ({new_n484_, new_n730_})
2'b11 : new_n4663_ = 1'b1;
default : new_n4663_ = 1'b0;
endcase
casez ({new_n96_, new_n451_})
2'b11 : new_n4664_ = 1'b1;
default : new_n4664_ = 1'b0;
endcase
casez ({new_n280_, new_n454_})
2'b11 : new_n4665_ = 1'b1;
default : new_n4665_ = 1'b0;
endcase
casez ({new_n80_, new_n457_})
2'b11 : new_n4666_ = 1'b1;
default : new_n4666_ = 1'b0;
endcase
casez ({y[2], new_n472_})
2'b01 : new_n4667_ = 1'b1;
default : new_n4667_ = 1'b0;
endcase
casez ({new_n103_, new_n473_})
2'b11 : new_n4668_ = 1'b1;
default : new_n4668_ = 1'b0;
endcase
casez ({new_n157_, new_n209_})
2'b11 : new_n4669_ = 1'b1;
default : new_n4669_ = 1'b0;
endcase
casez ({new_n646_, new_n1905_})
2'b00 : new_n4670_ = 1'b1;
default : new_n4670_ = 1'b0;
endcase
casez ({new_n1210_, new_n1907_})
2'b00 : new_n4671_ = 1'b1;
default : new_n4671_ = 1'b0;
endcase
casez ({new_n97_, new_n492_, new_n772_})
3'b10? : new_n4672_ = 1'b1;
3'b??1 : new_n4672_ = 1'b1;
default : new_n4672_ = 1'b0;
endcase
casez ({new_n463_, new_n777_})
2'b00 : new_n4673_ = 1'b1;
default : new_n4673_ = 1'b0;
endcase
casez ({new_n643_, new_n1927_})
2'b00 : new_n4674_ = 1'b1;
default : new_n4674_ = 1'b0;
endcase
casez ({new_n109_, new_n697_, new_n1927_})
3'b01? : new_n4675_ = 1'b1;
3'b??1 : new_n4675_ = 1'b1;
default : new_n4675_ = 1'b0;
endcase
casez ({new_n812_, new_n1928_})
2'b00 : new_n4676_ = 1'b1;
default : new_n4676_ = 1'b0;
endcase
casez ({new_n1710_, new_n1931_})
2'b10 : new_n4677_ = 1'b1;
default : new_n4677_ = 1'b0;
endcase
casez ({new_n289_, new_n490_})
2'b00 : new_n4678_ = 1'b1;
default : new_n4678_ = 1'b0;
endcase
casez ({new_n1484_, new_n1933_})
2'b00 : new_n4679_ = 1'b1;
default : new_n4679_ = 1'b0;
endcase
casez ({new_n1461_, new_n1934_})
2'b00 : new_n4680_ = 1'b1;
default : new_n4680_ = 1'b0;
endcase
casez ({new_n570_, new_n782_})
2'b00 : new_n4681_ = 1'b1;
default : new_n4681_ = 1'b0;
endcase
casez ({new_n94_, new_n720_, new_n109_, new_n1953_})
4'b10?? : new_n4682_ = 1'b1;
4'b??01 : new_n4682_ = 1'b1;
default : new_n4682_ = 1'b0;
endcase
casez ({new_n463_, new_n1164_})
2'b00 : new_n4683_ = 1'b1;
default : new_n4683_ = 1'b0;
endcase
casez ({new_n899_, new_n1164_})
2'b00 : new_n4684_ = 1'b1;
default : new_n4684_ = 1'b0;
endcase
casez ({new_n1034_, new_n1965_})
2'b01 : new_n4685_ = 1'b1;
default : new_n4685_ = 1'b0;
endcase
casez ({new_n188_, new_n787_})
2'b00 : new_n4686_ = 1'b1;
default : new_n4686_ = 1'b0;
endcase
casez ({new_n756_, new_n788_})
2'b00 : new_n4687_ = 1'b1;
default : new_n4687_ = 1'b0;
endcase
casez ({new_n645_, new_n788_})
2'b00 : new_n4688_ = 1'b1;
default : new_n4688_ = 1'b0;
endcase
casez ({new_n667_, new_n1969_})
2'b01 : new_n4689_ = 1'b1;
default : new_n4689_ = 1'b0;
endcase
casez ({new_n164_, new_n263_})
2'b00 : new_n4690_ = 1'b1;
default : new_n4690_ = 1'b0;
endcase
casez ({new_n412_, new_n503_})
2'b00 : new_n4691_ = 1'b1;
default : new_n4691_ = 1'b0;
endcase
casez ({new_n695_, new_n789_})
2'b00 : new_n4692_ = 1'b1;
default : new_n4692_ = 1'b0;
endcase
casez ({new_n1334_, new_n1980_})
2'b01 : new_n4693_ = 1'b1;
default : new_n4693_ = 1'b0;
endcase
casez ({new_n648_, new_n1176_})
2'b00 : new_n4694_ = 1'b1;
default : new_n4694_ = 1'b0;
endcase
casez ({new_n793_, new_n1997_})
2'b01 : new_n4695_ = 1'b1;
default : new_n4695_ = 1'b0;
endcase
casez ({new_n627_, new_n1998_})
2'b01 : new_n4696_ = 1'b1;
default : new_n4696_ = 1'b0;
endcase
casez ({new_n1866_, new_n2001_})
2'b01 : new_n4697_ = 1'b1;
default : new_n4697_ = 1'b0;
endcase
casez ({new_n520_, new_n1182_})
2'b00 : new_n4698_ = 1'b1;
default : new_n4698_ = 1'b0;
endcase
casez ({new_n197_, new_n797_})
2'b00 : new_n4699_ = 1'b1;
default : new_n4699_ = 1'b0;
endcase
casez ({new_n752_, new_n2024_})
2'b01 : new_n4700_ = 1'b1;
default : new_n4700_ = 1'b0;
endcase
casez ({new_n434_, new_n800_})
2'b00 : new_n4701_ = 1'b1;
default : new_n4701_ = 1'b0;
endcase
casez ({new_n455_, new_n520_})
2'b00 : new_n4702_ = 1'b1;
default : new_n4702_ = 1'b0;
endcase
casez ({new_n514_, new_n1199_})
2'b00 : new_n4703_ = 1'b1;
default : new_n4703_ = 1'b0;
endcase
casez ({new_n1018_, new_n1200_})
2'b00 : new_n4704_ = 1'b1;
default : new_n4704_ = 1'b0;
endcase
casez ({new_n856_, new_n1201_})
2'b00 : new_n4705_ = 1'b1;
default : new_n4705_ = 1'b0;
endcase
casez ({new_n723_, new_n1202_})
2'b00 : new_n4706_ = 1'b1;
default : new_n4706_ = 1'b0;
endcase
casez ({new_n1737_, new_n2058_})
2'b01 : new_n4707_ = 1'b1;
default : new_n4707_ = 1'b0;
endcase
casez ({new_n2051_, new_n2061_})
2'b11 : new_n4708_ = 1'b1;
default : new_n4708_ = 1'b0;
endcase
casez ({new_n1067_, new_n1204_})
2'b00 : new_n4709_ = 1'b1;
default : new_n4709_ = 1'b0;
endcase
casez ({new_n1874_, new_n2066_})
2'b01 : new_n4710_ = 1'b1;
default : new_n4710_ = 1'b0;
endcase
casez ({new_n496_, new_n2067_})
2'b01 : new_n4711_ = 1'b1;
default : new_n4711_ = 1'b0;
endcase
casez ({new_n1016_, new_n2069_})
2'b01 : new_n4712_ = 1'b1;
default : new_n4712_ = 1'b0;
endcase
casez ({new_n229_, new_n262_, new_n809_})
3'b11? : new_n4713_ = 1'b1;
3'b??1 : new_n4713_ = 1'b1;
default : new_n4713_ = 1'b0;
endcase
casez ({new_n1307_, new_n2072_})
2'b01 : new_n4714_ = 1'b1;
default : new_n4714_ = 1'b0;
endcase
casez ({new_n752_, new_n2081_})
2'b01 : new_n4715_ = 1'b1;
default : new_n4715_ = 1'b0;
endcase
casez ({new_n1113_, new_n2081_})
2'b01 : new_n4716_ = 1'b1;
default : new_n4716_ = 1'b0;
endcase
casez ({new_n245_, new_n533_})
2'b00 : new_n4717_ = 1'b1;
default : new_n4717_ = 1'b0;
endcase
casez ({new_n173_, new_n187_, new_n1210_})
3'b11? : new_n4718_ = 1'b1;
3'b??1 : new_n4718_ = 1'b1;
default : new_n4718_ = 1'b0;
endcase
casez ({new_n396_, new_n2091_})
2'b01 : new_n4719_ = 1'b1;
default : new_n4719_ = 1'b0;
endcase
casez ({new_n810_, new_n812_})
2'b00 : new_n4720_ = 1'b1;
default : new_n4720_ = 1'b0;
endcase
casez ({new_n2022_, new_n2094_})
2'b11 : new_n4721_ = 1'b1;
default : new_n4721_ = 1'b0;
endcase
casez ({new_n613_, new_n1212_})
2'b00 : new_n4722_ = 1'b1;
default : new_n4722_ = 1'b0;
endcase
casez ({new_n472_, new_n1212_})
2'b00 : new_n4723_ = 1'b1;
default : new_n4723_ = 1'b0;
endcase
casez ({new_n1066_, new_n1213_})
2'b00 : new_n4724_ = 1'b1;
default : new_n4724_ = 1'b0;
endcase
casez ({new_n974_, new_n2101_})
2'b01 : new_n4725_ = 1'b1;
default : new_n4725_ = 1'b0;
endcase
casez ({new_n1885_, new_n2103_})
2'b01 : new_n4726_ = 1'b1;
default : new_n4726_ = 1'b0;
endcase
casez ({new_n160_, new_n386_, new_n1214_})
3'b11? : new_n4727_ = 1'b1;
3'b??1 : new_n4727_ = 1'b1;
default : new_n4727_ = 1'b0;
endcase
casez ({new_n350_, new_n2104_})
2'b01 : new_n4728_ = 1'b1;
default : new_n4728_ = 1'b0;
endcase
casez ({new_n277_, new_n2105_})
2'b01 : new_n4729_ = 1'b1;
default : new_n4729_ = 1'b0;
endcase
casez ({new_n618_, new_n2107_})
2'b01 : new_n4730_ = 1'b1;
default : new_n4730_ = 1'b0;
endcase
casez ({new_n897_, new_n2107_})
2'b01 : new_n4731_ = 1'b1;
default : new_n4731_ = 1'b0;
endcase
casez ({new_n867_, new_n1214_})
2'b00 : new_n4732_ = 1'b1;
default : new_n4732_ = 1'b0;
endcase
casez ({new_n384_, new_n1215_})
2'b00 : new_n4733_ = 1'b1;
default : new_n4733_ = 1'b0;
endcase
casez ({new_n1203_, new_n2110_})
2'b00 : new_n4734_ = 1'b1;
default : new_n4734_ = 1'b0;
endcase
casez ({new_n1178_, new_n1215_})
2'b00 : new_n4735_ = 1'b1;
default : new_n4735_ = 1'b0;
endcase
casez ({new_n827_, new_n2110_})
2'b00 : new_n4736_ = 1'b1;
default : new_n4736_ = 1'b0;
endcase
casez ({new_n718_, new_n2111_})
2'b00 : new_n4737_ = 1'b1;
default : new_n4737_ = 1'b0;
endcase
casez ({new_n166_, new_n289_, new_n2112_})
3'b11? : new_n4738_ = 1'b1;
3'b??1 : new_n4738_ = 1'b1;
default : new_n4738_ = 1'b0;
endcase
casez ({new_n237_, new_n275_, new_n1216_})
3'b11? : new_n4739_ = 1'b1;
3'b??1 : new_n4739_ = 1'b1;
default : new_n4739_ = 1'b0;
endcase
casez ({new_n1594_, new_n2113_})
2'b00 : new_n4740_ = 1'b1;
default : new_n4740_ = 1'b0;
endcase
casez ({new_n814_, new_n816_})
2'b00 : new_n4741_ = 1'b1;
default : new_n4741_ = 1'b0;
endcase
casez ({new_n850_, new_n2116_})
2'b00 : new_n4742_ = 1'b1;
default : new_n4742_ = 1'b0;
endcase
casez ({new_n1109_, new_n1217_})
2'b00 : new_n4743_ = 1'b1;
default : new_n4743_ = 1'b0;
endcase
casez ({new_n1732_, new_n2117_})
2'b00 : new_n4744_ = 1'b1;
default : new_n4744_ = 1'b0;
endcase
casez ({new_n1152_, new_n2118_})
2'b00 : new_n4745_ = 1'b1;
default : new_n4745_ = 1'b0;
endcase
casez ({new_n948_, new_n2118_})
2'b00 : new_n4746_ = 1'b1;
default : new_n4746_ = 1'b0;
endcase
casez ({u[0], new_n494_, new_n2119_})
3'b01? : new_n4747_ = 1'b1;
3'b??1 : new_n4747_ = 1'b1;
default : new_n4747_ = 1'b0;
endcase
casez ({new_n1727_, new_n2119_})
2'b00 : new_n4748_ = 1'b1;
default : new_n4748_ = 1'b0;
endcase
casez ({new_n1203_, new_n2119_})
2'b00 : new_n4749_ = 1'b1;
default : new_n4749_ = 1'b0;
endcase
casez ({new_n1223_, new_n2120_})
2'b00 : new_n4750_ = 1'b1;
default : new_n4750_ = 1'b0;
endcase
casez ({new_n1287_, new_n2120_})
2'b00 : new_n4751_ = 1'b1;
default : new_n4751_ = 1'b0;
endcase
casez ({new_n445_, new_n936_, new_n1219_})
3'b10? : new_n4752_ = 1'b1;
3'b??1 : new_n4752_ = 1'b1;
default : new_n4752_ = 1'b0;
endcase
casez ({new_n1227_, new_n2121_})
2'b00 : new_n4753_ = 1'b1;
default : new_n4753_ = 1'b0;
endcase
casez ({new_n1131_, new_n2121_})
2'b00 : new_n4754_ = 1'b1;
default : new_n4754_ = 1'b0;
endcase
casez ({new_n1592_, new_n2122_})
2'b00 : new_n4755_ = 1'b1;
default : new_n4755_ = 1'b0;
endcase
casez ({new_n1375_, new_n2122_})
2'b00 : new_n4756_ = 1'b1;
default : new_n4756_ = 1'b0;
endcase
casez ({new_n980_, new_n2122_})
2'b00 : new_n4757_ = 1'b1;
default : new_n4757_ = 1'b0;
endcase
casez ({new_n1065_, new_n2122_})
2'b00 : new_n4758_ = 1'b1;
default : new_n4758_ = 1'b0;
endcase
casez ({new_n647_, new_n1221_})
2'b00 : new_n4759_ = 1'b1;
default : new_n4759_ = 1'b0;
endcase
casez ({new_n718_, new_n2125_})
2'b00 : new_n4760_ = 1'b1;
default : new_n4760_ = 1'b0;
endcase
casez ({new_n570_, new_n1221_})
2'b00 : new_n4761_ = 1'b1;
default : new_n4761_ = 1'b0;
endcase
casez ({new_n1105_, new_n2128_})
2'b00 : new_n4762_ = 1'b1;
default : new_n4762_ = 1'b0;
endcase
casez ({new_n738_, new_n2128_})
2'b00 : new_n4763_ = 1'b1;
default : new_n4763_ = 1'b0;
endcase
casez ({new_n904_, new_n2129_})
2'b00 : new_n4764_ = 1'b1;
default : new_n4764_ = 1'b0;
endcase
casez ({new_n663_, new_n1223_})
2'b00 : new_n4765_ = 1'b1;
default : new_n4765_ = 1'b0;
endcase
casez ({new_n908_, new_n2130_})
2'b00 : new_n4766_ = 1'b1;
default : new_n4766_ = 1'b0;
endcase
casez ({new_n92_, new_n2130_, new_n193_, new_n228_})
4'b01?? : new_n4767_ = 1'b1;
4'b??11 : new_n4767_ = 1'b1;
default : new_n4767_ = 1'b0;
endcase
casez ({new_n983_, new_n2131_})
2'b00 : new_n4768_ = 1'b1;
default : new_n4768_ = 1'b0;
endcase
casez ({new_n756_, new_n2131_})
2'b00 : new_n4769_ = 1'b1;
default : new_n4769_ = 1'b0;
endcase
casez ({new_n581_, new_n2132_})
2'b00 : new_n4770_ = 1'b1;
default : new_n4770_ = 1'b0;
endcase
casez ({new_n955_, new_n1224_})
2'b00 : new_n4771_ = 1'b1;
default : new_n4771_ = 1'b0;
endcase
casez ({new_n1225_, new_n2133_})
2'b00 : new_n4772_ = 1'b1;
default : new_n4772_ = 1'b0;
endcase
casez ({new_n1346_, new_n2134_})
2'b00 : new_n4773_ = 1'b1;
default : new_n4773_ = 1'b0;
endcase
casez ({new_n1223_, new_n2134_})
2'b00 : new_n4774_ = 1'b1;
default : new_n4774_ = 1'b0;
endcase
casez ({new_n121_, new_n317_, new_n1226_})
3'b11? : new_n4775_ = 1'b1;
3'b??1 : new_n4775_ = 1'b1;
default : new_n4775_ = 1'b0;
endcase
casez ({new_n186_, new_n254_, new_n2136_})
3'b11? : new_n4776_ = 1'b1;
3'b??1 : new_n4776_ = 1'b1;
default : new_n4776_ = 1'b0;
endcase
casez ({new_n212_, new_n385_, new_n2137_})
3'b11? : new_n4777_ = 1'b1;
3'b??1 : new_n4777_ = 1'b1;
default : new_n4777_ = 1'b0;
endcase
casez ({new_n1058_, new_n2138_})
2'b00 : new_n4778_ = 1'b1;
default : new_n4778_ = 1'b0;
endcase
casez ({new_n1376_, new_n2138_})
2'b00 : new_n4779_ = 1'b1;
default : new_n4779_ = 1'b0;
endcase
casez ({new_n1213_, new_n2139_})
2'b00 : new_n4780_ = 1'b1;
default : new_n4780_ = 1'b0;
endcase
casez ({new_n639_, new_n1227_})
2'b00 : new_n4781_ = 1'b1;
default : new_n4781_ = 1'b0;
endcase
casez ({new_n1216_, new_n2140_})
2'b00 : new_n4782_ = 1'b1;
default : new_n4782_ = 1'b0;
endcase
casez ({new_n2132_, new_n2140_})
2'b00 : new_n4783_ = 1'b1;
default : new_n4783_ = 1'b0;
endcase
casez ({new_n118_, new_n239_, new_n828_})
3'b11? : new_n4784_ = 1'b1;
3'b??1 : new_n4784_ = 1'b1;
default : new_n4784_ = 1'b0;
endcase
casez ({new_n402_, new_n1227_})
2'b00 : new_n4785_ = 1'b1;
default : new_n4785_ = 1'b0;
endcase
casez ({new_n84_, new_n829_, new_n637_})
3'b11? : new_n4786_ = 1'b1;
3'b??1 : new_n4786_ = 1'b1;
default : new_n4786_ = 1'b0;
endcase
casez ({new_n724_, new_n2141_})
2'b00 : new_n4787_ = 1'b1;
default : new_n4787_ = 1'b0;
endcase
casez ({new_n1157_, new_n2142_})
2'b00 : new_n4788_ = 1'b1;
default : new_n4788_ = 1'b0;
endcase
casez ({new_n540_, new_n544_})
2'b00 : new_n4789_ = 1'b1;
default : new_n4789_ = 1'b0;
endcase
casez ({new_n754_, new_n830_})
2'b00 : new_n4790_ = 1'b1;
default : new_n4790_ = 1'b0;
endcase
casez ({new_n1377_, new_n2143_})
2'b00 : new_n4791_ = 1'b1;
default : new_n4791_ = 1'b0;
endcase
casez ({new_n1739_, new_n2143_})
2'b00 : new_n4792_ = 1'b1;
default : new_n4792_ = 1'b0;
endcase
casez ({new_n1481_, new_n2144_})
2'b00 : new_n4793_ = 1'b1;
default : new_n4793_ = 1'b0;
endcase
casez ({new_n199_, new_n260_, new_n544_})
3'b11? : new_n4794_ = 1'b1;
3'b??1 : new_n4794_ = 1'b1;
default : new_n4794_ = 1'b0;
endcase
casez ({new_n1904_, new_n2145_})
2'b00 : new_n4795_ = 1'b1;
default : new_n4795_ = 1'b0;
endcase
casez ({new_n755_, new_n834_})
2'b00 : new_n4796_ = 1'b1;
default : new_n4796_ = 1'b0;
endcase
casez ({new_n899_, new_n2148_})
2'b00 : new_n4797_ = 1'b1;
default : new_n4797_ = 1'b0;
endcase
casez ({v[1], new_n2150_, new_n89_, new_n340_})
4'b01?? : new_n4798_ = 1'b1;
4'b??11 : new_n4798_ = 1'b1;
default : new_n4798_ = 1'b0;
endcase
casez ({new_n603_, new_n2150_})
2'b00 : new_n4799_ = 1'b1;
default : new_n4799_ = 1'b0;
endcase
casez ({new_n5435_, new_n287_, new_n329_})
3'b1?? : new_n4800_ = 1'b1;
3'b?11 : new_n4800_ = 1'b1;
default : new_n4800_ = 1'b0;
endcase
casez ({new_n510_, new_n836_})
2'b00 : new_n4801_ = 1'b1;
default : new_n4801_ = 1'b0;
endcase
casez ({new_n826_, new_n2152_})
2'b00 : new_n4802_ = 1'b1;
default : new_n4802_ = 1'b0;
endcase
casez ({new_n625_, new_n2152_})
2'b00 : new_n4803_ = 1'b1;
default : new_n4803_ = 1'b0;
endcase
casez ({new_n667_, new_n2152_})
2'b00 : new_n4804_ = 1'b1;
default : new_n4804_ = 1'b0;
endcase
casez ({new_n816_, new_n2153_})
2'b00 : new_n4805_ = 1'b1;
default : new_n4805_ = 1'b0;
endcase
casez ({new_n2115_, new_n2155_})
2'b00 : new_n4806_ = 1'b1;
default : new_n4806_ = 1'b0;
endcase
casez ({new_n104_, new_n2156_, new_n1717_})
3'b01? : new_n4807_ = 1'b1;
3'b??1 : new_n4807_ = 1'b1;
default : new_n4807_ = 1'b0;
endcase
casez ({new_n1466_, new_n2160_})
2'b00 : new_n4808_ = 1'b1;
default : new_n4808_ = 1'b0;
endcase
casez ({new_n666_, new_n2160_})
2'b00 : new_n4809_ = 1'b1;
default : new_n4809_ = 1'b0;
endcase
casez ({new_n1041_, new_n2161_})
2'b00 : new_n4810_ = 1'b1;
default : new_n4810_ = 1'b0;
endcase
casez ({new_n552_, new_n845_})
2'b00 : new_n4811_ = 1'b1;
default : new_n4811_ = 1'b0;
endcase
casez ({new_n214_, new_n422_, new_n850_})
3'b11? : new_n4812_ = 1'b1;
3'b??1 : new_n4812_ = 1'b1;
default : new_n4812_ = 1'b0;
endcase
casez ({new_n520_, new_n851_})
2'b00 : new_n4813_ = 1'b1;
default : new_n4813_ = 1'b0;
endcase
casez ({new_n848_, new_n852_})
2'b00 : new_n4814_ = 1'b1;
default : new_n4814_ = 1'b0;
endcase
casez ({new_n367_, new_n561_})
2'b00 : new_n4815_ = 1'b1;
default : new_n4815_ = 1'b0;
endcase
casez ({new_n717_, new_n1270_})
2'b00 : new_n4816_ = 1'b1;
default : new_n4816_ = 1'b0;
endcase
casez ({new_n848_, new_n1273_})
2'b00 : new_n4817_ = 1'b1;
default : new_n4817_ = 1'b0;
endcase
casez ({new_n658_, new_n1273_})
2'b00 : new_n4818_ = 1'b1;
default : new_n4818_ = 1'b0;
endcase
casez ({new_n1141_, new_n1277_})
2'b00 : new_n4819_ = 1'b1;
default : new_n4819_ = 1'b0;
endcase
casez ({new_n482_, new_n1280_})
2'b00 : new_n4820_ = 1'b1;
default : new_n4820_ = 1'b0;
endcase
casez ({new_n494_, new_n1283_})
2'b00 : new_n4821_ = 1'b1;
default : new_n4821_ = 1'b0;
endcase
casez ({new_n900_, new_n1285_})
2'b00 : new_n4822_ = 1'b1;
default : new_n4822_ = 1'b0;
endcase
casez ({new_n566_, new_n1285_})
2'b00 : new_n4823_ = 1'b1;
default : new_n4823_ = 1'b0;
endcase
casez ({new_n144_, new_n369_, new_n1293_})
3'b11? : new_n4824_ = 1'b1;
3'b??1 : new_n4824_ = 1'b1;
default : new_n4824_ = 1'b0;
endcase
casez ({v[1], new_n318_, new_n1294_})
3'b11? : new_n4825_ = 1'b1;
3'b??1 : new_n4825_ = 1'b1;
default : new_n4825_ = 1'b0;
endcase
casez ({new_n600_, new_n1295_})
2'b00 : new_n4826_ = 1'b1;
default : new_n4826_ = 1'b0;
endcase
casez ({new_n985_, new_n1300_})
2'b00 : new_n4827_ = 1'b1;
default : new_n4827_ = 1'b0;
endcase
casez ({new_n154_, new_n598_, new_n1301_})
3'b11? : new_n4828_ = 1'b1;
3'b??1 : new_n4828_ = 1'b1;
default : new_n4828_ = 1'b0;
endcase
casez ({new_n189_, new_n1305_, new_n625_})
3'b10? : new_n4829_ = 1'b1;
3'b??1 : new_n4829_ = 1'b1;
default : new_n4829_ = 1'b0;
endcase
casez ({new_n109_, new_n199_, new_n569_})
3'b01? : new_n4830_ = 1'b1;
3'b??1 : new_n4830_ = 1'b1;
default : new_n4830_ = 1'b0;
endcase
casez ({new_n625_, new_n1312_})
2'b00 : new_n4831_ = 1'b1;
default : new_n4831_ = 1'b0;
endcase
casez ({new_n391_, new_n1320_})
2'b00 : new_n4832_ = 1'b1;
default : new_n4832_ = 1'b0;
endcase
casez ({new_n1055_, new_n1320_})
2'b00 : new_n4833_ = 1'b1;
default : new_n4833_ = 1'b0;
endcase
casez ({new_n350_, new_n572_})
2'b00 : new_n4834_ = 1'b1;
default : new_n4834_ = 1'b0;
endcase
casez ({new_n513_, new_n1323_})
2'b00 : new_n4835_ = 1'b1;
default : new_n4835_ = 1'b0;
endcase
casez ({x[0], new_n407_, new_n1324_})
3'b01? : new_n4836_ = 1'b1;
3'b??1 : new_n4836_ = 1'b1;
default : new_n4836_ = 1'b0;
endcase
casez ({new_n643_, new_n1328_})
2'b00 : new_n4837_ = 1'b1;
default : new_n4837_ = 1'b0;
endcase
casez ({new_n238_, new_n576_})
2'b00 : new_n4838_ = 1'b1;
default : new_n4838_ = 1'b0;
endcase
casez ({new_n277_, new_n297_})
2'b00 : new_n4839_ = 1'b1;
default : new_n4839_ = 1'b0;
endcase
casez ({new_n5453_, new_n1332_})
2'b1? : new_n4840_ = 1'b1;
2'b?1 : new_n4840_ = 1'b1;
default : new_n4840_ = 1'b0;
endcase
casez ({new_n109_, new_n405_, new_n1332_})
3'b01? : new_n4841_ = 1'b1;
3'b??1 : new_n4841_ = 1'b1;
default : new_n4841_ = 1'b0;
endcase
casez ({new_n1070_, new_n1333_})
2'b00 : new_n4842_ = 1'b1;
default : new_n4842_ = 1'b0;
endcase
casez ({new_n1108_, new_n1334_})
2'b00 : new_n4843_ = 1'b1;
default : new_n4843_ = 1'b0;
endcase
casez ({new_n1295_, new_n1336_})
2'b00 : new_n4844_ = 1'b1;
default : new_n4844_ = 1'b0;
endcase
casez ({new_n814_, new_n1339_})
2'b00 : new_n4845_ = 1'b1;
default : new_n4845_ = 1'b0;
endcase
casez ({new_n1203_, new_n1340_})
2'b00 : new_n4846_ = 1'b1;
default : new_n4846_ = 1'b0;
endcase
casez ({new_n613_, new_n1340_})
2'b00 : new_n4847_ = 1'b1;
default : new_n4847_ = 1'b0;
endcase
casez ({x[1], new_n987_, new_n1343_})
3'b11? : new_n4848_ = 1'b1;
3'b??1 : new_n4848_ = 1'b1;
default : new_n4848_ = 1'b0;
endcase
casez ({new_n561_, new_n1345_})
2'b00 : new_n4849_ = 1'b1;
default : new_n4849_ = 1'b0;
endcase
casez ({new_n649_, new_n1349_})
2'b00 : new_n4850_ = 1'b1;
default : new_n4850_ = 1'b0;
endcase
casez ({new_n440_, new_n1354_})
2'b00 : new_n4851_ = 1'b1;
default : new_n4851_ = 1'b0;
endcase
casez ({new_n836_, new_n1356_})
2'b00 : new_n4852_ = 1'b1;
default : new_n4852_ = 1'b0;
endcase
casez ({new_n98_, new_n240_, new_n897_})
3'b11? : new_n4853_ = 1'b1;
3'b??1 : new_n4853_ = 1'b1;
default : new_n4853_ = 1'b0;
endcase
casez ({new_n978_, new_n1358_})
2'b00 : new_n4854_ = 1'b1;
default : new_n4854_ = 1'b0;
endcase
casez ({new_n717_, new_n897_})
2'b00 : new_n4855_ = 1'b1;
default : new_n4855_ = 1'b0;
endcase
casez ({new_n242_, new_n488_, new_n901_})
3'b11? : new_n4856_ = 1'b1;
3'b??1 : new_n4856_ = 1'b1;
default : new_n4856_ = 1'b0;
endcase
casez ({new_n610_, new_n902_})
2'b00 : new_n4857_ = 1'b1;
default : new_n4857_ = 1'b0;
endcase
casez ({new_n169_, new_n220_, new_n903_})
3'b11? : new_n4858_ = 1'b1;
3'b??1 : new_n4858_ = 1'b1;
default : new_n4858_ = 1'b0;
endcase
casez ({new_n577_, new_n903_})
2'b00 : new_n4859_ = 1'b1;
default : new_n4859_ = 1'b0;
endcase
casez ({new_n376_, new_n1373_})
2'b00 : new_n4860_ = 1'b1;
default : new_n4860_ = 1'b0;
endcase
casez ({new_n723_, new_n904_})
2'b00 : new_n4861_ = 1'b1;
default : new_n4861_ = 1'b0;
endcase
casez ({new_n402_, new_n905_})
2'b00 : new_n4862_ = 1'b1;
default : new_n4862_ = 1'b0;
endcase
casez ({new_n463_, new_n905_})
2'b00 : new_n4863_ = 1'b1;
default : new_n4863_ = 1'b0;
endcase
casez ({new_n544_, new_n905_})
2'b00 : new_n4864_ = 1'b1;
default : new_n4864_ = 1'b0;
endcase
casez ({new_n727_, new_n1378_})
2'b00 : new_n4865_ = 1'b1;
default : new_n4865_ = 1'b0;
endcase
casez ({new_n984_, new_n1379_})
2'b00 : new_n4866_ = 1'b1;
default : new_n4866_ = 1'b0;
endcase
casez ({new_n611_, new_n1380_})
2'b00 : new_n4867_ = 1'b1;
default : new_n4867_ = 1'b0;
endcase
casez ({new_n813_, new_n1380_})
2'b00 : new_n4868_ = 1'b1;
default : new_n4868_ = 1'b0;
endcase
casez ({new_n724_, new_n908_})
2'b00 : new_n4869_ = 1'b1;
default : new_n4869_ = 1'b0;
endcase
casez ({new_n647_, new_n909_})
2'b00 : new_n4870_ = 1'b1;
default : new_n4870_ = 1'b0;
endcase
casez ({new_n577_, new_n910_})
2'b00 : new_n4871_ = 1'b1;
default : new_n4871_ = 1'b0;
endcase
casez ({new_n534_, new_n1387_})
2'b00 : new_n4872_ = 1'b1;
default : new_n4872_ = 1'b0;
endcase
casez ({new_n1322_, new_n1391_})
2'b00 : new_n4873_ = 1'b1;
default : new_n4873_ = 1'b0;
endcase
casez ({new_n572_, new_n1393_})
2'b00 : new_n4874_ = 1'b1;
default : new_n4874_ = 1'b0;
endcase
casez ({new_n158_, new_n2524_, new_n168_, new_n1261_})
4'b11?? : new_n4875_ = 1'b1;
4'b??10 : new_n4875_ = 1'b1;
default : new_n4875_ = 1'b0;
endcase
casez ({new_n255_, new_n2539_, new_n976_})
3'b10? : new_n4876_ = 1'b1;
3'b??1 : new_n4876_ = 1'b1;
default : new_n4876_ = 1'b0;
endcase
casez ({new_n131_, new_n2541_, new_n1479_})
3'b10? : new_n4877_ = 1'b1;
3'b??1 : new_n4877_ = 1'b1;
default : new_n4877_ = 1'b0;
endcase
casez ({new_n181_, new_n1703_, new_n236_, new_n2553_})
4'b00?? : new_n4878_ = 1'b1;
4'b??11 : new_n4878_ = 1'b1;
default : new_n4878_ = 1'b0;
endcase
casez ({new_n2064_, new_n2554_})
2'b10 : new_n4879_ = 1'b1;
default : new_n4879_ = 1'b0;
endcase
casez ({new_n434_, new_n1394_})
2'b00 : new_n4880_ = 1'b1;
default : new_n4880_ = 1'b0;
endcase
casez ({new_n1214_, new_n2563_})
2'b00 : new_n4881_ = 1'b1;
default : new_n4881_ = 1'b0;
endcase
casez ({new_n191_, new_n469_, new_n613_})
3'b11? : new_n4882_ = 1'b1;
3'b??1 : new_n4882_ = 1'b1;
default : new_n4882_ = 1'b0;
endcase
casez ({new_n1330_, new_n1399_})
2'b00 : new_n4883_ = 1'b1;
default : new_n4883_ = 1'b0;
endcase
casez ({new_n188_, new_n1400_})
2'b00 : new_n4884_ = 1'b1;
default : new_n4884_ = 1'b0;
endcase
casez ({new_n645_, new_n2572_})
2'b00 : new_n4885_ = 1'b1;
default : new_n4885_ = 1'b0;
endcase
casez ({new_n613_, new_n2577_})
2'b00 : new_n4886_ = 1'b1;
default : new_n4886_ = 1'b0;
endcase
casez ({new_n1488_, new_n2580_})
2'b00 : new_n4887_ = 1'b1;
default : new_n4887_ = 1'b0;
endcase
casez ({new_n2124_, new_n2581_})
2'b00 : new_n4888_ = 1'b1;
default : new_n4888_ = 1'b0;
endcase
casez ({new_n263_, new_n2583_})
2'b00 : new_n4889_ = 1'b1;
default : new_n4889_ = 1'b0;
endcase
casez ({new_n816_, new_n2587_})
2'b00 : new_n4890_ = 1'b1;
default : new_n4890_ = 1'b0;
endcase
casez ({new_n373_, new_n1409_})
2'b01 : new_n4891_ = 1'b1;
default : new_n4891_ = 1'b0;
endcase
casez ({new_n646_, new_n2590_})
2'b00 : new_n4892_ = 1'b1;
default : new_n4892_ = 1'b0;
endcase
casez ({new_n484_, new_n1409_})
2'b01 : new_n4893_ = 1'b1;
default : new_n4893_ = 1'b0;
endcase
casez ({new_n842_, new_n1413_})
2'b01 : new_n4894_ = 1'b1;
default : new_n4894_ = 1'b0;
endcase
casez ({new_n296_, new_n618_})
2'b00 : new_n4895_ = 1'b1;
default : new_n4895_ = 1'b0;
endcase
casez ({new_n177_, new_n927_, new_n725_})
3'b11? : new_n4896_ = 1'b1;
3'b??1 : new_n4896_ = 1'b1;
default : new_n4896_ = 1'b0;
endcase
casez ({new_n113_, new_n932_, new_n904_})
3'b11? : new_n4897_ = 1'b1;
3'b??1 : new_n4897_ = 1'b1;
default : new_n4897_ = 1'b0;
endcase
casez ({new_n1205_, new_n2620_})
2'b00 : new_n4898_ = 1'b1;
default : new_n4898_ = 1'b0;
endcase
casez ({new_n1056_, new_n1438_})
2'b01 : new_n4899_ = 1'b1;
default : new_n4899_ = 1'b0;
endcase
casez ({new_n612_, new_n623_})
2'b00 : new_n4900_ = 1'b1;
default : new_n4900_ = 1'b0;
endcase
casez ({new_n368_, new_n623_})
2'b00 : new_n4901_ = 1'b1;
default : new_n4901_ = 1'b0;
endcase
casez ({new_n835_, new_n2634_})
2'b00 : new_n4902_ = 1'b1;
default : new_n4902_ = 1'b0;
endcase
casez ({new_n195_, new_n1447_})
2'b01 : new_n4903_ = 1'b1;
default : new_n4903_ = 1'b0;
endcase
casez ({new_n1393_, new_n1447_})
2'b01 : new_n4904_ = 1'b1;
default : new_n4904_ = 1'b0;
endcase
casez ({new_n613_, new_n2637_})
2'b00 : new_n4905_ = 1'b1;
default : new_n4905_ = 1'b0;
endcase
casez ({new_n644_, new_n2643_})
2'b00 : new_n4906_ = 1'b1;
default : new_n4906_ = 1'b0;
endcase
casez ({new_n96_, new_n2646_, new_n625_})
3'b01? : new_n4907_ = 1'b1;
3'b??1 : new_n4907_ = 1'b1;
default : new_n4907_ = 1'b0;
endcase
casez ({new_n1038_, new_n1455_})
2'b01 : new_n4908_ = 1'b1;
default : new_n4908_ = 1'b0;
endcase
casez ({new_n2127_, new_n2649_})
2'b00 : new_n4909_ = 1'b1;
default : new_n4909_ = 1'b0;
endcase
casez ({new_n1200_, new_n2651_})
2'b00 : new_n4910_ = 1'b1;
default : new_n4910_ = 1'b0;
endcase
casez ({new_n637_, new_n1457_})
2'b00 : new_n4911_ = 1'b1;
default : new_n4911_ = 1'b0;
endcase
casez ({new_n204_, new_n240_, new_n1458_})
3'b11? : new_n4912_ = 1'b1;
3'b??1 : new_n4912_ = 1'b1;
default : new_n4912_ = 1'b0;
endcase
casez ({new_n96_, new_n668_, new_n1459_})
3'b11? : new_n4913_ = 1'b1;
3'b??1 : new_n4913_ = 1'b1;
default : new_n4913_ = 1'b0;
endcase
casez ({new_n1055_, new_n1459_})
2'b00 : new_n4914_ = 1'b1;
default : new_n4914_ = 1'b0;
endcase
casez ({new_n1734_, new_n2661_})
2'b00 : new_n4915_ = 1'b1;
default : new_n4915_ = 1'b0;
endcase
casez ({new_n463_, new_n944_})
2'b00 : new_n4916_ = 1'b1;
default : new_n4916_ = 1'b0;
endcase
casez ({new_n1123_, new_n1460_})
2'b00 : new_n4917_ = 1'b1;
default : new_n4917_ = 1'b0;
endcase
casez ({new_n645_, new_n2665_})
2'b00 : new_n4918_ = 1'b1;
default : new_n4918_ = 1'b0;
endcase
casez ({new_n568_, new_n945_})
2'b00 : new_n4919_ = 1'b1;
default : new_n4919_ = 1'b0;
endcase
casez ({new_n1204_, new_n2670_})
2'b00 : new_n4920_ = 1'b1;
default : new_n4920_ = 1'b0;
endcase
casez ({new_n1721_, new_n2670_})
2'b00 : new_n4921_ = 1'b1;
default : new_n4921_ = 1'b0;
endcase
casez ({new_n215_, new_n332_, new_n1462_})
3'b11? : new_n4922_ = 1'b1;
3'b??1 : new_n4922_ = 1'b1;
default : new_n4922_ = 1'b0;
endcase
casez ({new_n322_, new_n336_})
2'b00 : new_n4923_ = 1'b1;
default : new_n4923_ = 1'b0;
endcase
casez ({new_n1731_, new_n2673_})
2'b00 : new_n4924_ = 1'b1;
default : new_n4924_ = 1'b0;
endcase
casez ({new_n245_, new_n1464_})
2'b00 : new_n4925_ = 1'b1;
default : new_n4925_ = 1'b0;
endcase
casez ({new_n462_, new_n2676_})
2'b00 : new_n4926_ = 1'b1;
default : new_n4926_ = 1'b0;
endcase
casez ({new_n900_, new_n1465_})
2'b00 : new_n4927_ = 1'b1;
default : new_n4927_ = 1'b0;
endcase
casez ({new_n84_, new_n713_, new_n1466_})
3'b11? : new_n4928_ = 1'b1;
3'b??1 : new_n4928_ = 1'b1;
default : new_n4928_ = 1'b0;
endcase
casez ({new_n721_, new_n1467_})
2'b10 : new_n4929_ = 1'b1;
default : new_n4929_ = 1'b0;
endcase
casez ({new_n1216_, new_n1467_})
2'b00 : new_n4930_ = 1'b1;
default : new_n4930_ = 1'b0;
endcase
casez ({new_n2131_, new_n2696_})
2'b00 : new_n4931_ = 1'b1;
default : new_n4931_ = 1'b0;
endcase
casez ({new_n1462_, new_n2696_})
2'b00 : new_n4932_ = 1'b1;
default : new_n4932_ = 1'b0;
endcase
casez ({new_n624_, new_n2696_})
2'b00 : new_n4933_ = 1'b1;
default : new_n4933_ = 1'b0;
endcase
casez ({new_n535_, new_n1469_})
2'b00 : new_n4934_ = 1'b1;
default : new_n4934_ = 1'b0;
endcase
casez ({new_n723_, new_n951_})
2'b00 : new_n4935_ = 1'b1;
default : new_n4935_ = 1'b0;
endcase
casez ({new_n968_, new_n2712_})
2'b10 : new_n4936_ = 1'b1;
default : new_n4936_ = 1'b0;
endcase
casez ({new_n867_, new_n1474_})
2'b00 : new_n4937_ = 1'b1;
default : new_n4937_ = 1'b0;
endcase
casez ({new_n1206_, new_n2715_})
2'b00 : new_n4938_ = 1'b1;
default : new_n4938_ = 1'b0;
endcase
casez ({new_n1207_, new_n1475_})
2'b00 : new_n4939_ = 1'b1;
default : new_n4939_ = 1'b0;
endcase
casez ({new_n1433_, new_n2720_})
2'b10 : new_n4940_ = 1'b1;
default : new_n4940_ = 1'b0;
endcase
casez ({new_n976_, new_n1476_})
2'b00 : new_n4941_ = 1'b1;
default : new_n4941_ = 1'b0;
endcase
casez ({new_n1748_, new_n2721_})
2'b00 : new_n4942_ = 1'b1;
default : new_n4942_ = 1'b0;
endcase
casez ({new_n1302_, new_n2722_})
2'b00 : new_n4943_ = 1'b1;
default : new_n4943_ = 1'b0;
endcase
casez ({new_n611_, new_n1476_})
2'b00 : new_n4944_ = 1'b1;
default : new_n4944_ = 1'b0;
endcase
casez ({new_n642_, new_n1477_})
2'b00 : new_n4945_ = 1'b1;
default : new_n4945_ = 1'b0;
endcase
casez ({new_n2151_, new_n2725_})
2'b00 : new_n4946_ = 1'b1;
default : new_n4946_ = 1'b0;
endcase
casez ({new_n854_, new_n1477_})
2'b00 : new_n4947_ = 1'b1;
default : new_n4947_ = 1'b0;
endcase
casez ({new_n646_, new_n1478_})
2'b00 : new_n4948_ = 1'b1;
default : new_n4948_ = 1'b0;
endcase
casez ({new_n390_, new_n925_, new_n1480_})
3'b10? : new_n4949_ = 1'b1;
3'b??1 : new_n4949_ = 1'b1;
default : new_n4949_ = 1'b0;
endcase
casez ({new_n642_, new_n2740_})
2'b00 : new_n4950_ = 1'b1;
default : new_n4950_ = 1'b0;
endcase
casez ({new_n434_, new_n2741_})
2'b00 : new_n4951_ = 1'b1;
default : new_n4951_ = 1'b0;
endcase
casez ({new_n1213_, new_n1483_})
2'b00 : new_n4952_ = 1'b1;
default : new_n4952_ = 1'b0;
endcase
casez ({new_n88_, new_n639_, new_n624_})
3'b01? : new_n4953_ = 1'b1;
3'b??1 : new_n4953_ = 1'b1;
default : new_n4953_ = 1'b0;
endcase
casez ({new_n544_, new_n2751_})
2'b00 : new_n4954_ = 1'b1;
default : new_n4954_ = 1'b0;
endcase
casez ({new_n677_, new_n1484_})
2'b00 : new_n4955_ = 1'b1;
default : new_n4955_ = 1'b0;
endcase
casez ({new_n569_, new_n639_})
2'b00 : new_n4956_ = 1'b1;
default : new_n4956_ = 1'b0;
endcase
casez ({new_n845_, new_n2760_})
2'b00 : new_n4957_ = 1'b1;
default : new_n4957_ = 1'b0;
endcase
casez ({new_n800_, new_n1486_})
2'b00 : new_n4958_ = 1'b1;
default : new_n4958_ = 1'b0;
endcase
casez ({new_n2072_, new_n2761_})
2'b10 : new_n4959_ = 1'b1;
default : new_n4959_ = 1'b0;
endcase
casez ({new_n176_, new_n219_, new_n1487_})
3'b11? : new_n4960_ = 1'b1;
3'b??1 : new_n4960_ = 1'b1;
default : new_n4960_ = 1'b0;
endcase
casez ({new_n1223_, new_n1488_})
2'b00 : new_n4961_ = 1'b1;
default : new_n4961_ = 1'b0;
endcase
casez ({new_n477_, new_n1488_})
2'b00 : new_n4962_ = 1'b1;
default : new_n4962_ = 1'b0;
endcase
casez ({new_n1466_, new_n2766_})
2'b00 : new_n4963_ = 1'b1;
default : new_n4963_ = 1'b0;
endcase
casez ({new_n745_, new_n1488_})
2'b00 : new_n4964_ = 1'b1;
default : new_n4964_ = 1'b0;
endcase
casez ({new_n96_, new_n2769_, new_n1480_})
3'b01? : new_n4965_ = 1'b1;
3'b??1 : new_n4965_ = 1'b1;
default : new_n4965_ = 1'b0;
endcase
casez ({new_n695_, new_n962_})
2'b00 : new_n4966_ = 1'b1;
default : new_n4966_ = 1'b0;
endcase
casez ({new_n1329_, new_n2776_})
2'b00 : new_n4967_ = 1'b1;
default : new_n4967_ = 1'b0;
endcase
casez ({new_n860_, new_n1491_})
2'b00 : new_n4968_ = 1'b1;
default : new_n4968_ = 1'b0;
endcase
casez ({new_n89_, new_n620_, new_n1492_})
3'b01? : new_n4969_ = 1'b1;
3'b??1 : new_n4969_ = 1'b1;
default : new_n4969_ = 1'b0;
endcase
casez ({new_n1314_, new_n2779_})
2'b00 : new_n4970_ = 1'b1;
default : new_n4970_ = 1'b0;
endcase
casez ({new_n755_, new_n963_})
2'b00 : new_n4971_ = 1'b1;
default : new_n4971_ = 1'b0;
endcase
casez ({new_n148_, new_n2782_, new_n610_})
3'b10? : new_n4972_ = 1'b1;
3'b??1 : new_n4972_ = 1'b1;
default : new_n4972_ = 1'b0;
endcase
casez ({new_n97_, new_n1132_, new_n166_, new_n2785_})
4'b11?? : new_n4973_ = 1'b1;
4'b??10 : new_n4973_ = 1'b1;
default : new_n4973_ = 1'b0;
endcase
casez ({new_n440_, new_n1492_})
2'b00 : new_n4974_ = 1'b1;
default : new_n4974_ = 1'b0;
endcase
casez ({new_n141_, new_n2789_, new_n308_, new_n712_})
4'b11?? : new_n4975_ = 1'b1;
4'b??11 : new_n4975_ = 1'b1;
default : new_n4975_ = 1'b0;
endcase
casez ({new_n1651_, new_n2789_})
2'b00 : new_n4976_ = 1'b1;
default : new_n4976_ = 1'b0;
endcase
casez ({new_n1746_, new_n2790_})
2'b00 : new_n4977_ = 1'b1;
default : new_n4977_ = 1'b0;
endcase
casez ({new_n904_, new_n2790_})
2'b00 : new_n4978_ = 1'b1;
default : new_n4978_ = 1'b0;
endcase
casez ({new_n631_, new_n2791_})
2'b00 : new_n4979_ = 1'b1;
default : new_n4979_ = 1'b0;
endcase
casez ({new_n1714_, new_n2792_})
2'b00 : new_n4980_ = 1'b1;
default : new_n4980_ = 1'b0;
endcase
casez ({new_n1862_, new_n2792_})
2'b00 : new_n4981_ = 1'b1;
default : new_n4981_ = 1'b0;
endcase
casez ({new_n976_, new_n2794_})
2'b00 : new_n4982_ = 1'b1;
default : new_n4982_ = 1'b0;
endcase
casez ({new_n506_, new_n644_})
2'b00 : new_n4983_ = 1'b1;
default : new_n4983_ = 1'b0;
endcase
casez ({new_n83_, new_n1721_, new_n2798_})
3'b01? : new_n4984_ = 1'b1;
3'b??1 : new_n4984_ = 1'b1;
default : new_n4984_ = 1'b0;
endcase
casez ({new_n1728_, new_n2799_})
2'b00 : new_n4985_ = 1'b1;
default : new_n4985_ = 1'b0;
endcase
casez ({new_n148_, new_n966_, new_n241_, new_n393_})
4'b10?? : new_n4986_ = 1'b1;
4'b??10 : new_n4986_ = 1'b1;
default : new_n4986_ = 1'b0;
endcase
casez ({new_n1036_, new_n2802_})
2'b00 : new_n4987_ = 1'b1;
default : new_n4987_ = 1'b0;
endcase
casez ({new_n201_, new_n338_, new_n1498_})
3'b11? : new_n4988_ = 1'b1;
3'b??1 : new_n4988_ = 1'b1;
default : new_n4988_ = 1'b0;
endcase
casez ({new_n455_, new_n971_})
2'b01 : new_n4989_ = 1'b1;
default : new_n4989_ = 1'b0;
endcase
casez ({new_n678_, new_n2803_})
2'b00 : new_n4990_ = 1'b1;
default : new_n4990_ = 1'b0;
endcase
casez ({new_n1131_, new_n1498_})
2'b00 : new_n4991_ = 1'b1;
default : new_n4991_ = 1'b0;
endcase
casez ({new_n251_, new_n261_, new_n2803_})
3'b11? : new_n4992_ = 1'b1;
3'b??1 : new_n4992_ = 1'b1;
default : new_n4992_ = 1'b0;
endcase
casez ({new_n164_, new_n971_, new_n306_, new_n441_})
4'b10?? : new_n4993_ = 1'b1;
4'b??11 : new_n4993_ = 1'b1;
default : new_n4993_ = 1'b0;
endcase
casez ({new_n865_, new_n2808_})
2'b00 : new_n4994_ = 1'b1;
default : new_n4994_ = 1'b0;
endcase
casez ({new_n1164_, new_n1500_})
2'b00 : new_n4995_ = 1'b1;
default : new_n4995_ = 1'b0;
endcase
casez ({new_n2141_, new_n2808_})
2'b00 : new_n4996_ = 1'b1;
default : new_n4996_ = 1'b0;
endcase
casez ({new_n899_, new_n2809_})
2'b00 : new_n4997_ = 1'b1;
default : new_n4997_ = 1'b0;
endcase
casez ({new_n755_, new_n1501_})
2'b00 : new_n4998_ = 1'b1;
default : new_n4998_ = 1'b0;
endcase
casez ({new_n746_, new_n2810_})
2'b00 : new_n4999_ = 1'b1;
default : new_n4999_ = 1'b0;
endcase
casez ({new_n1067_, new_n2810_})
2'b00 : new_n5000_ = 1'b1;
default : new_n5000_ = 1'b0;
endcase
casez ({new_n1342_, new_n2811_})
2'b00 : new_n5001_ = 1'b1;
default : new_n5001_ = 1'b0;
endcase
casez ({new_n1359_, new_n2811_})
2'b00 : new_n5002_ = 1'b1;
default : new_n5002_ = 1'b0;
endcase
casez ({new_n981_, new_n2812_})
2'b00 : new_n5003_ = 1'b1;
default : new_n5003_ = 1'b0;
endcase
casez ({new_n2724_, new_n2812_})
2'b00 : new_n5004_ = 1'b1;
default : new_n5004_ = 1'b0;
endcase
casez ({new_n1899_, new_n2813_})
2'b00 : new_n5005_ = 1'b1;
default : new_n5005_ = 1'b0;
endcase
casez ({new_n657_, new_n973_})
2'b00 : new_n5006_ = 1'b1;
default : new_n5006_ = 1'b0;
endcase
casez ({new_n899_, new_n1502_})
2'b00 : new_n5007_ = 1'b1;
default : new_n5007_ = 1'b0;
endcase
casez ({new_n223_, new_n493_, new_n1502_})
3'b11? : new_n5008_ = 1'b1;
3'b??1 : new_n5008_ = 1'b1;
default : new_n5008_ = 1'b0;
endcase
casez ({new_n463_, new_n2814_})
2'b00 : new_n5009_ = 1'b1;
default : new_n5009_ = 1'b0;
endcase
casez ({new_n947_, new_n974_})
2'b00 : new_n5010_ = 1'b1;
default : new_n5010_ = 1'b0;
endcase
casez ({new_n951_, new_n2815_})
2'b00 : new_n5011_ = 1'b1;
default : new_n5011_ = 1'b0;
endcase
casez ({new_n151_, new_n228_, new_n2815_})
3'b11? : new_n5012_ = 1'b1;
3'b??1 : new_n5012_ = 1'b1;
default : new_n5012_ = 1'b0;
endcase
casez ({new_n973_, new_n2817_})
2'b00 : new_n5013_ = 1'b1;
default : new_n5013_ = 1'b0;
endcase
casez ({new_n2121_, new_n2818_})
2'b00 : new_n5014_ = 1'b1;
default : new_n5014_ = 1'b0;
endcase
casez ({new_n1227_, new_n1505_})
2'b00 : new_n5015_ = 1'b1;
default : new_n5015_ = 1'b0;
endcase
casez ({new_n659_, new_n716_, new_n2821_})
3'b01? : new_n5016_ = 1'b1;
3'b??1 : new_n5016_ = 1'b1;
default : new_n5016_ = 1'b0;
endcase
casez ({new_n905_, new_n1505_})
2'b00 : new_n5017_ = 1'b1;
default : new_n5017_ = 1'b0;
endcase
casez ({new_n1027_, new_n2822_})
2'b00 : new_n5018_ = 1'b1;
default : new_n5018_ = 1'b0;
endcase
casez ({new_n1028_, new_n2824_})
2'b00 : new_n5019_ = 1'b1;
default : new_n5019_ = 1'b0;
endcase
casez ({new_n755_, new_n2824_})
2'b00 : new_n5020_ = 1'b1;
default : new_n5020_ = 1'b0;
endcase
casez ({new_n463_, new_n2825_})
2'b00 : new_n5021_ = 1'b1;
default : new_n5021_ = 1'b0;
endcase
casez ({new_n2129_, new_n2826_})
2'b00 : new_n5022_ = 1'b1;
default : new_n5022_ = 1'b0;
endcase
casez ({new_n1472_, new_n2827_})
2'b00 : new_n5023_ = 1'b1;
default : new_n5023_ = 1'b0;
endcase
casez ({new_n426_, new_n1539_, new_n2827_})
3'b11? : new_n5024_ = 1'b1;
3'b??1 : new_n5024_ = 1'b1;
default : new_n5024_ = 1'b0;
endcase
casez ({new_n1469_, new_n2828_})
2'b00 : new_n5025_ = 1'b1;
default : new_n5025_ = 1'b0;
endcase
casez ({new_n269_, new_n355_})
2'b00 : new_n5026_ = 1'b1;
default : new_n5026_ = 1'b0;
endcase
casez ({new_n740_, new_n2831_})
2'b00 : new_n5027_ = 1'b1;
default : new_n5027_ = 1'b0;
endcase
casez ({new_n416_, new_n2835_})
2'b00 : new_n5028_ = 1'b1;
default : new_n5028_ = 1'b0;
endcase
casez ({new_n954_, new_n977_})
2'b00 : new_n5029_ = 1'b1;
default : new_n5029_ = 1'b0;
endcase
casez ({new_n480_, new_n2547_, new_n2841_})
3'b10? : new_n5030_ = 1'b1;
3'b??1 : new_n5030_ = 1'b1;
default : new_n5030_ = 1'b0;
endcase
casez ({new_n81_, new_n483_, new_n2841_})
3'b01? : new_n5031_ = 1'b1;
3'b??1 : new_n5031_ = 1'b1;
default : new_n5031_ = 1'b0;
endcase
casez ({new_n789_, new_n2842_})
2'b00 : new_n5032_ = 1'b1;
default : new_n5032_ = 1'b0;
endcase
casez ({new_n430_, new_n633_, new_n2845_})
3'b11? : new_n5033_ = 1'b1;
3'b??1 : new_n5033_ = 1'b1;
default : new_n5033_ = 1'b0;
endcase
casez ({new_n325_, new_n648_})
2'b00 : new_n5034_ = 1'b1;
default : new_n5034_ = 1'b0;
endcase
casez ({new_n1141_, new_n2848_})
2'b00 : new_n5035_ = 1'b1;
default : new_n5035_ = 1'b0;
endcase
casez ({new_n720_, new_n2848_})
2'b10 : new_n5036_ = 1'b1;
default : new_n5036_ = 1'b0;
endcase
casez ({new_n942_, new_n981_})
2'b00 : new_n5037_ = 1'b1;
default : new_n5037_ = 1'b0;
endcase
casez ({new_n378_, new_n982_})
2'b00 : new_n5038_ = 1'b1;
default : new_n5038_ = 1'b0;
endcase
casez ({new_n646_, new_n983_})
2'b00 : new_n5039_ = 1'b1;
default : new_n5039_ = 1'b0;
endcase
casez ({new_n666_, new_n983_})
2'b00 : new_n5040_ = 1'b1;
default : new_n5040_ = 1'b0;
endcase
casez ({new_n908_, new_n986_})
2'b00 : new_n5041_ = 1'b1;
default : new_n5041_ = 1'b0;
endcase
casez ({new_n1162_, new_n1553_})
2'b00 : new_n5042_ = 1'b1;
default : new_n5042_ = 1'b0;
endcase
casez ({new_n164_, new_n338_, new_n988_})
3'b11? : new_n5043_ = 1'b1;
3'b??1 : new_n5043_ = 1'b1;
default : new_n5043_ = 1'b0;
endcase
casez ({new_n726_, new_n1560_})
2'b00 : new_n5044_ = 1'b1;
default : new_n5044_ = 1'b0;
endcase
casez ({new_n83_, new_n350_, new_n665_})
3'b11? : new_n5045_ = 1'b1;
3'b??1 : new_n5045_ = 1'b1;
default : new_n5045_ = 1'b0;
endcase
casez ({new_n981_, new_n1561_})
2'b00 : new_n5046_ = 1'b1;
default : new_n5046_ = 1'b0;
endcase
casez ({new_n770_, new_n2952_})
2'b00 : new_n5047_ = 1'b1;
default : new_n5047_ = 1'b0;
endcase
casez ({new_n1313_, new_n1563_})
2'b00 : new_n5048_ = 1'b1;
default : new_n5048_ = 1'b0;
endcase
casez ({new_n1307_, new_n1565_})
2'b00 : new_n5049_ = 1'b1;
default : new_n5049_ = 1'b0;
endcase
casez ({new_n795_, new_n995_})
2'b00 : new_n5050_ = 1'b1;
default : new_n5050_ = 1'b0;
endcase
casez ({new_n932_, new_n1567_})
2'b00 : new_n5051_ = 1'b1;
default : new_n5051_ = 1'b0;
endcase
casez ({new_n524_, new_n2982_})
2'b00 : new_n5052_ = 1'b1;
default : new_n5052_ = 1'b0;
endcase
casez ({new_n1920_, new_n2985_})
2'b00 : new_n5053_ = 1'b1;
default : new_n5053_ = 1'b0;
endcase
casez ({new_n1737_, new_n2987_})
2'b00 : new_n5054_ = 1'b1;
default : new_n5054_ = 1'b0;
endcase
casez ({new_n901_, new_n2994_})
2'b00 : new_n5055_ = 1'b1;
default : new_n5055_ = 1'b0;
endcase
casez ({new_n947_, new_n2999_})
2'b00 : new_n5056_ = 1'b1;
default : new_n5056_ = 1'b0;
endcase
casez ({x[1], new_n347_, new_n3002_})
3'b11? : new_n5057_ = 1'b1;
3'b??1 : new_n5057_ = 1'b1;
default : new_n5057_ = 1'b0;
endcase
casez ({u[0], new_n435_, new_n3003_})
3'b01? : new_n5058_ = 1'b1;
3'b??1 : new_n5058_ = 1'b1;
default : new_n5058_ = 1'b0;
endcase
casez ({new_n2832_, new_n3008_})
2'b00 : new_n5059_ = 1'b1;
default : new_n5059_ = 1'b0;
endcase
casez ({new_n2751_, new_n3011_})
2'b00 : new_n5060_ = 1'b1;
default : new_n5060_ = 1'b0;
endcase
casez ({new_n867_, new_n3015_})
2'b00 : new_n5061_ = 1'b1;
default : new_n5061_ = 1'b0;
endcase
casez ({new_n698_, new_n1003_})
2'b00 : new_n5062_ = 1'b1;
default : new_n5062_ = 1'b0;
endcase
casez ({new_n84_, new_n221_, new_n373_})
3'b11? : new_n5063_ = 1'b1;
3'b??1 : new_n5063_ = 1'b1;
default : new_n5063_ = 1'b0;
endcase
casez ({new_n1364_, new_n3021_})
2'b00 : new_n5064_ = 1'b1;
default : new_n5064_ = 1'b0;
endcase
casez ({new_n949_, new_n3033_})
2'b00 : new_n5065_ = 1'b1;
default : new_n5065_ = 1'b0;
endcase
casez ({new_n647_, new_n1004_})
2'b00 : new_n5066_ = 1'b1;
default : new_n5066_ = 1'b0;
endcase
casez ({new_n255_, new_n363_, new_n3035_})
3'b11? : new_n5067_ = 1'b1;
3'b??1 : new_n5067_ = 1'b1;
default : new_n5067_ = 1'b0;
endcase
casez ({new_n2951_, new_n2967_, new_n3036_})
3'b11? : new_n5068_ = 1'b1;
3'b??1 : new_n5068_ = 1'b1;
default : new_n5068_ = 1'b0;
endcase
casez ({new_n583_, new_n3038_})
2'b00 : new_n5069_ = 1'b1;
default : new_n5069_ = 1'b0;
endcase
casez ({new_n85_, new_n1796_, new_n3044_})
3'b11? : new_n5070_ = 1'b1;
3'b??1 : new_n5070_ = 1'b1;
default : new_n5070_ = 1'b0;
endcase
casez ({new_n1964_, new_n3053_})
2'b00 : new_n5071_ = 1'b1;
default : new_n5071_ = 1'b0;
endcase
casez ({new_n1106_, new_n3055_})
2'b00 : new_n5072_ = 1'b1;
default : new_n5072_ = 1'b0;
endcase
casez ({new_n121_, new_n493_, new_n3056_})
3'b11? : new_n5073_ = 1'b1;
3'b??1 : new_n5073_ = 1'b1;
default : new_n5073_ = 1'b0;
endcase
casez ({new_n2161_, new_n3071_})
2'b00 : new_n5074_ = 1'b1;
default : new_n5074_ = 1'b0;
endcase
casez ({new_n1736_, new_n3072_})
2'b00 : new_n5075_ = 1'b1;
default : new_n5075_ = 1'b0;
endcase
casez ({new_n1716_, new_n3076_})
2'b00 : new_n5076_ = 1'b1;
default : new_n5076_ = 1'b0;
endcase
casez ({new_n1502_, new_n3078_})
2'b00 : new_n5077_ = 1'b1;
default : new_n5077_ = 1'b0;
endcase
casez ({new_n1891_, new_n3082_})
2'b00 : new_n5078_ = 1'b1;
default : new_n5078_ = 1'b0;
endcase
casez ({new_n1105_, new_n3086_})
2'b00 : new_n5079_ = 1'b1;
default : new_n5079_ = 1'b0;
endcase
casez ({new_n236_, new_n3089_})
2'b00 : new_n5080_ = 1'b1;
default : new_n5080_ = 1'b0;
endcase
casez ({new_n1623_, new_n3094_})
2'b00 : new_n5081_ = 1'b1;
default : new_n5081_ = 1'b0;
endcase
casez ({new_n1159_, new_n3096_})
2'b00 : new_n5082_ = 1'b1;
default : new_n5082_ = 1'b0;
endcase
casez ({new_n177_, new_n244_, new_n3097_})
3'b11? : new_n5083_ = 1'b1;
3'b??1 : new_n5083_ = 1'b1;
default : new_n5083_ = 1'b0;
endcase
casez ({new_n1827_, new_n3106_})
2'b00 : new_n5084_ = 1'b1;
default : new_n5084_ = 1'b0;
endcase
casez ({new_n1287_, new_n1585_})
2'b00 : new_n5085_ = 1'b1;
default : new_n5085_ = 1'b0;
endcase
casez ({new_n1045_, new_n3108_})
2'b00 : new_n5086_ = 1'b1;
default : new_n5086_ = 1'b0;
endcase
casez ({new_n2564_, new_n3114_})
2'b00 : new_n5087_ = 1'b1;
default : new_n5087_ = 1'b0;
endcase
casez ({new_n2111_, new_n3115_})
2'b00 : new_n5088_ = 1'b1;
default : new_n5088_ = 1'b0;
endcase
casez ({new_n527_, new_n3116_})
2'b00 : new_n5089_ = 1'b1;
default : new_n5089_ = 1'b0;
endcase
casez ({new_n2661_, new_n3120_})
2'b00 : new_n5090_ = 1'b1;
default : new_n5090_ = 1'b0;
endcase
casez ({new_n1606_, new_n3124_})
2'b00 : new_n5091_ = 1'b1;
default : new_n5091_ = 1'b0;
endcase
casez ({new_n1394_, new_n3126_})
2'b00 : new_n5092_ = 1'b1;
default : new_n5092_ = 1'b0;
endcase
casez ({new_n627_, new_n3130_})
2'b01 : new_n5093_ = 1'b1;
default : new_n5093_ = 1'b0;
endcase
casez ({new_n373_, new_n3142_})
2'b00 : new_n5094_ = 1'b1;
default : new_n5094_ = 1'b0;
endcase
casez ({new_n105_, new_n3145_})
2'b00 : new_n5095_ = 1'b1;
default : new_n5095_ = 1'b0;
endcase
casez ({new_n1357_, new_n3146_})
2'b00 : new_n5096_ = 1'b1;
default : new_n5096_ = 1'b0;
endcase
casez ({new_n739_, new_n3149_})
2'b00 : new_n5097_ = 1'b1;
default : new_n5097_ = 1'b0;
endcase
casez ({new_n84_, new_n734_, new_n3156_})
3'b11? : new_n5098_ = 1'b1;
3'b??1 : new_n5098_ = 1'b1;
default : new_n5098_ = 1'b0;
endcase
casez ({new_n1391_, new_n3158_})
2'b00 : new_n5099_ = 1'b1;
default : new_n5099_ = 1'b0;
endcase
casez ({new_n1218_, new_n3166_})
2'b00 : new_n5100_ = 1'b1;
default : new_n5100_ = 1'b0;
endcase
casez ({new_n1922_, new_n3167_})
2'b00 : new_n5101_ = 1'b1;
default : new_n5101_ = 1'b0;
endcase
casez ({new_n646_, new_n1015_})
2'b00 : new_n5102_ = 1'b1;
default : new_n5102_ = 1'b0;
endcase
casez ({new_n974_, new_n1015_})
2'b00 : new_n5103_ = 1'b1;
default : new_n5103_ = 1'b0;
endcase
casez ({new_n1465_, new_n3172_})
2'b00 : new_n5104_ = 1'b1;
default : new_n5104_ = 1'b0;
endcase
casez ({new_n172_, new_n1091_, new_n3174_})
3'b10? : new_n5105_ = 1'b1;
3'b??1 : new_n5105_ = 1'b1;
default : new_n5105_ = 1'b0;
endcase
casez ({new_n2622_, new_n3183_})
2'b00 : new_n5106_ = 1'b1;
default : new_n5106_ = 1'b0;
endcase
casez ({new_n1283_, new_n3184_})
2'b00 : new_n5107_ = 1'b1;
default : new_n5107_ = 1'b0;
endcase
casez ({new_n1299_, new_n3185_})
2'b00 : new_n5108_ = 1'b1;
default : new_n5108_ = 1'b0;
endcase
casez ({new_n1859_, new_n3186_})
2'b00 : new_n5109_ = 1'b1;
default : new_n5109_ = 1'b0;
endcase
casez ({new_n983_, new_n1596_})
2'b00 : new_n5110_ = 1'b1;
default : new_n5110_ = 1'b0;
endcase
casez ({new_n2925_, new_n3189_})
2'b00 : new_n5111_ = 1'b1;
default : new_n5111_ = 1'b0;
endcase
casez ({new_n498_, new_n3193_})
2'b00 : new_n5112_ = 1'b1;
default : new_n5112_ = 1'b0;
endcase
casez ({new_n1293_, new_n3194_})
2'b00 : new_n5113_ = 1'b1;
default : new_n5113_ = 1'b0;
endcase
casez ({new_n958_, new_n3195_})
2'b00 : new_n5114_ = 1'b1;
default : new_n5114_ = 1'b0;
endcase
casez ({new_n624_, new_n3198_})
2'b00 : new_n5115_ = 1'b1;
default : new_n5115_ = 1'b0;
endcase
casez ({new_n1392_, new_n3199_})
2'b00 : new_n5116_ = 1'b1;
default : new_n5116_ = 1'b0;
endcase
casez ({new_n1309_, new_n1598_})
2'b00 : new_n5117_ = 1'b1;
default : new_n5117_ = 1'b0;
endcase
casez ({new_n645_, new_n1599_})
2'b00 : new_n5118_ = 1'b1;
default : new_n5118_ = 1'b0;
endcase
casez ({new_n807_, new_n3212_})
2'b00 : new_n5119_ = 1'b1;
default : new_n5119_ = 1'b0;
endcase
casez ({new_n1392_, new_n3214_})
2'b00 : new_n5120_ = 1'b1;
default : new_n5120_ = 1'b0;
endcase
casez ({new_n1914_, new_n3230_})
2'b00 : new_n5121_ = 1'b1;
default : new_n5121_ = 1'b0;
endcase
casez ({new_n791_, new_n3231_})
2'b00 : new_n5122_ = 1'b1;
default : new_n5122_ = 1'b0;
endcase
casez ({new_n1292_, new_n3237_})
2'b00 : new_n5123_ = 1'b1;
default : new_n5123_ = 1'b0;
endcase
casez ({new_n2599_, new_n3245_})
2'b00 : new_n5124_ = 1'b1;
default : new_n5124_ = 1'b0;
endcase
casez ({new_n678_, new_n3246_})
2'b00 : new_n5125_ = 1'b1;
default : new_n5125_ = 1'b0;
endcase
casez ({new_n708_, new_n1020_})
2'b00 : new_n5126_ = 1'b1;
default : new_n5126_ = 1'b0;
endcase
casez ({new_n1623_, new_n3256_})
2'b00 : new_n5127_ = 1'b1;
default : new_n5127_ = 1'b0;
endcase
casez ({new_n1489_, new_n3261_})
2'b00 : new_n5128_ = 1'b1;
default : new_n5128_ = 1'b0;
endcase
casez ({new_n1738_, new_n3267_})
2'b00 : new_n5129_ = 1'b1;
default : new_n5129_ = 1'b0;
endcase
casez ({new_n665_, new_n3268_})
2'b00 : new_n5130_ = 1'b1;
default : new_n5130_ = 1'b0;
endcase
casez ({new_n131_, new_n2530_, new_n3269_})
3'b10? : new_n5131_ = 1'b1;
3'b??1 : new_n5131_ = 1'b1;
default : new_n5131_ = 1'b0;
endcase
casez ({new_n1467_, new_n3270_})
2'b00 : new_n5132_ = 1'b1;
default : new_n5132_ = 1'b0;
endcase
casez ({new_n663_, new_n1608_})
2'b00 : new_n5133_ = 1'b1;
default : new_n5133_ = 1'b0;
endcase
casez ({new_n975_, new_n3274_})
2'b00 : new_n5134_ = 1'b1;
default : new_n5134_ = 1'b0;
endcase
casez ({new_n580_, new_n3277_})
2'b00 : new_n5135_ = 1'b1;
default : new_n5135_ = 1'b0;
endcase
casez ({new_n561_, new_n1609_})
2'b00 : new_n5136_ = 1'b1;
default : new_n5136_ = 1'b0;
endcase
casez ({new_n1611_, new_n3292_})
2'b00 : new_n5137_ = 1'b1;
default : new_n5137_ = 1'b0;
endcase
casez ({u[1], new_n290_, new_n3305_})
3'b11? : new_n5138_ = 1'b1;
3'b??1 : new_n5138_ = 1'b1;
default : new_n5138_ = 1'b0;
endcase
casez ({new_n240_, new_n719_, new_n3306_})
3'b11? : new_n5139_ = 1'b1;
3'b??1 : new_n5139_ = 1'b1;
default : new_n5139_ = 1'b0;
endcase
casez ({new_n1059_, new_n3307_})
2'b00 : new_n5140_ = 1'b1;
default : new_n5140_ = 1'b0;
endcase
casez ({new_n506_, new_n1612_})
2'b00 : new_n5141_ = 1'b1;
default : new_n5141_ = 1'b0;
endcase
casez ({new_n1632_, new_n3309_})
2'b00 : new_n5142_ = 1'b1;
default : new_n5142_ = 1'b0;
endcase
casez ({new_n373_, new_n3313_})
2'b00 : new_n5143_ = 1'b1;
default : new_n5143_ = 1'b0;
endcase
casez ({new_n506_, new_n3319_})
2'b00 : new_n5144_ = 1'b1;
default : new_n5144_ = 1'b0;
endcase
casez ({new_n646_, new_n3321_})
2'b00 : new_n5145_ = 1'b1;
default : new_n5145_ = 1'b0;
endcase
casez ({new_n756_, new_n1027_})
2'b00 : new_n5146_ = 1'b1;
default : new_n5146_ = 1'b0;
endcase
casez ({new_n1745_, new_n3324_})
2'b00 : new_n5147_ = 1'b1;
default : new_n5147_ = 1'b0;
endcase
casez ({new_n1738_, new_n3330_})
2'b00 : new_n5148_ = 1'b1;
default : new_n5148_ = 1'b0;
endcase
casez ({new_n1465_, new_n3337_})
2'b00 : new_n5149_ = 1'b1;
default : new_n5149_ = 1'b0;
endcase
casez ({new_n1457_, new_n3358_})
2'b00 : new_n5150_ = 1'b1;
default : new_n5150_ = 1'b0;
endcase
casez ({new_n373_, new_n1622_})
2'b00 : new_n5151_ = 1'b1;
default : new_n5151_ = 1'b0;
endcase
casez ({new_n825_, new_n1623_})
2'b00 : new_n5152_ = 1'b1;
default : new_n5152_ = 1'b0;
endcase
casez ({new_n2022_, new_n3366_})
2'b10 : new_n5153_ = 1'b1;
default : new_n5153_ = 1'b0;
endcase
casez ({new_n666_, new_n1624_})
2'b00 : new_n5154_ = 1'b1;
default : new_n5154_ = 1'b0;
endcase
casez ({new_n646_, new_n3385_})
2'b00 : new_n5155_ = 1'b1;
default : new_n5155_ = 1'b0;
endcase
casez ({new_n3023_, new_n3386_})
2'b00 : new_n5156_ = 1'b1;
default : new_n5156_ = 1'b0;
endcase
casez ({new_n909_, new_n3387_})
2'b00 : new_n5157_ = 1'b1;
default : new_n5157_ = 1'b0;
endcase
casez ({new_n1496_, new_n3393_})
2'b00 : new_n5158_ = 1'b1;
default : new_n5158_ = 1'b0;
endcase
casez ({new_n645_, new_n3406_})
2'b00 : new_n5159_ = 1'b1;
default : new_n5159_ = 1'b0;
endcase
casez ({new_n2152_, new_n3409_})
2'b00 : new_n5160_ = 1'b1;
default : new_n5160_ = 1'b0;
endcase
casez ({new_n131_, new_n179_, new_n696_})
3'b11? : new_n5161_ = 1'b1;
3'b??1 : new_n5161_ = 1'b1;
default : new_n5161_ = 1'b0;
endcase
casez ({new_n841_, new_n3432_})
2'b00 : new_n5162_ = 1'b1;
default : new_n5162_ = 1'b0;
endcase
casez ({new_n910_, new_n1037_})
2'b00 : new_n5163_ = 1'b1;
default : new_n5163_ = 1'b0;
endcase
casez ({new_n1054_, new_n3449_})
2'b00 : new_n5164_ = 1'b1;
default : new_n5164_ = 1'b0;
endcase
casez ({new_n1999_, new_n3450_})
2'b10 : new_n5165_ = 1'b1;
default : new_n5165_ = 1'b0;
endcase
casez ({new_n467_, new_n1038_})
2'b00 : new_n5166_ = 1'b1;
default : new_n5166_ = 1'b0;
endcase
casez ({new_n533_, new_n1038_})
2'b00 : new_n5167_ = 1'b1;
default : new_n5167_ = 1'b0;
endcase
casez ({new_n1734_, new_n3479_})
2'b00 : new_n5168_ = 1'b1;
default : new_n5168_ = 1'b0;
endcase
casez ({new_n1465_, new_n3488_})
2'b00 : new_n5169_ = 1'b1;
default : new_n5169_ = 1'b0;
endcase
casez ({new_n837_, new_n3490_})
2'b00 : new_n5170_ = 1'b1;
default : new_n5170_ = 1'b0;
endcase
casez ({new_n807_, new_n1041_})
2'b00 : new_n5171_ = 1'b1;
default : new_n5171_ = 1'b0;
endcase
casez ({new_n1221_, new_n3508_})
2'b00 : new_n5172_ = 1'b1;
default : new_n5172_ = 1'b0;
endcase
casez ({new_n1449_, new_n1648_})
2'b10 : new_n5173_ = 1'b1;
default : new_n5173_ = 1'b0;
endcase
casez ({x[1], new_n1650_, new_n561_})
3'b01? : new_n5174_ = 1'b1;
3'b??1 : new_n5174_ = 1'b1;
default : new_n5174_ = 1'b0;
endcase
casez ({new_n984_, new_n3542_})
2'b00 : new_n5175_ = 1'b1;
default : new_n5175_ = 1'b0;
endcase
casez ({new_n979_, new_n3548_})
2'b00 : new_n5176_ = 1'b1;
default : new_n5176_ = 1'b0;
endcase
casez ({new_n648_, new_n3559_})
2'b00 : new_n5177_ = 1'b1;
default : new_n5177_ = 1'b0;
endcase
casez ({new_n1423_, new_n3574_})
2'b10 : new_n5178_ = 1'b1;
default : new_n5178_ = 1'b0;
endcase
casez ({new_n515_, new_n3578_})
2'b00 : new_n5179_ = 1'b1;
default : new_n5179_ = 1'b0;
endcase
casez ({new_n97_, new_n706_, new_n373_})
3'b11? : new_n5180_ = 1'b1;
3'b??1 : new_n5180_ = 1'b1;
default : new_n5180_ = 1'b0;
endcase
casez ({new_n979_, new_n3593_})
2'b00 : new_n5181_ = 1'b1;
default : new_n5181_ = 1'b0;
endcase
casez ({new_n464_, new_n710_})
2'b00 : new_n5182_ = 1'b1;
default : new_n5182_ = 1'b0;
endcase
casez ({new_n1213_, new_n3604_})
2'b00 : new_n5183_ = 1'b1;
default : new_n5183_ = 1'b0;
endcase
casez ({new_n1722_, new_n3607_})
2'b00 : new_n5184_ = 1'b1;
default : new_n5184_ = 1'b0;
endcase
casez ({new_n538_, new_n3610_})
2'b01 : new_n5185_ = 1'b1;
default : new_n5185_ = 1'b0;
endcase
casez ({new_n516_, new_n710_})
2'b00 : new_n5186_ = 1'b1;
default : new_n5186_ = 1'b0;
endcase
casez ({new_n469_, new_n481_, new_n1054_})
3'b11? : new_n5187_ = 1'b1;
3'b??1 : new_n5187_ = 1'b1;
default : new_n5187_ = 1'b0;
endcase
casez ({new_n1225_, new_n3621_})
2'b01 : new_n5188_ = 1'b1;
default : new_n5188_ = 1'b0;
endcase
casez ({new_n2596_, new_n3624_})
2'b01 : new_n5189_ = 1'b1;
default : new_n5189_ = 1'b0;
endcase
casez ({new_n959_, new_n1054_})
2'b00 : new_n5190_ = 1'b1;
default : new_n5190_ = 1'b0;
endcase
casez ({new_n1011_, new_n1054_})
2'b00 : new_n5191_ = 1'b1;
default : new_n5191_ = 1'b0;
endcase
casez ({new_n512_, new_n3628_})
2'b01 : new_n5192_ = 1'b1;
default : new_n5192_ = 1'b0;
endcase
casez ({new_n1279_, new_n3629_})
2'b01 : new_n5193_ = 1'b1;
default : new_n5193_ = 1'b0;
endcase
casez ({u[2], new_n2540_, new_n3630_})
3'b00? : new_n5194_ = 1'b1;
3'b??0 : new_n5194_ = 1'b1;
default : new_n5194_ = 1'b0;
endcase
casez ({new_n2707_, new_n3631_})
2'b01 : new_n5195_ = 1'b1;
default : new_n5195_ = 1'b0;
endcase
casez ({new_n3077_, new_n3633_})
2'b01 : new_n5196_ = 1'b1;
default : new_n5196_ = 1'b0;
endcase
casez ({new_n2051_, new_n3639_})
2'b11 : new_n5197_ = 1'b1;
default : new_n5197_ = 1'b0;
endcase
casez ({new_n2663_, new_n3644_})
2'b01 : new_n5198_ = 1'b1;
default : new_n5198_ = 1'b0;
endcase
casez ({new_n754_, new_n1055_})
2'b00 : new_n5199_ = 1'b1;
default : new_n5199_ = 1'b0;
endcase
casez ({new_n1381_, new_n3649_})
2'b01 : new_n5200_ = 1'b1;
default : new_n5200_ = 1'b0;
endcase
casez ({new_n92_, new_n269_, new_n1055_})
3'b11? : new_n5201_ = 1'b1;
3'b??1 : new_n5201_ = 1'b1;
default : new_n5201_ = 1'b0;
endcase
casez ({new_n2578_, new_n3663_})
2'b01 : new_n5202_ = 1'b1;
default : new_n5202_ = 1'b0;
endcase
casez ({new_n1059_, new_n3680_})
2'b01 : new_n5203_ = 1'b1;
default : new_n5203_ = 1'b0;
endcase
casez ({new_n1316_, new_n3695_})
2'b01 : new_n5204_ = 1'b1;
default : new_n5204_ = 1'b0;
endcase
casez ({new_n1635_, new_n3703_})
2'b01 : new_n5205_ = 1'b1;
default : new_n5205_ = 1'b0;
endcase
casez ({new_n455_, new_n3706_})
2'b01 : new_n5206_ = 1'b1;
default : new_n5206_ = 1'b0;
endcase
casez ({new_n104_, new_n123_, new_n1712_})
3'b11? : new_n5207_ = 1'b1;
3'b??1 : new_n5207_ = 1'b1;
default : new_n5207_ = 1'b0;
endcase
casez ({x[2], new_n372_, new_n1712_})
3'b01? : new_n5208_ = 1'b1;
3'b??1 : new_n5208_ = 1'b1;
default : new_n5208_ = 1'b0;
endcase
casez ({new_n1633_, new_n3717_})
2'b01 : new_n5209_ = 1'b1;
default : new_n5209_ = 1'b0;
endcase
casez ({new_n907_, new_n1712_})
2'b00 : new_n5210_ = 1'b1;
default : new_n5210_ = 1'b0;
endcase
casez ({new_n1724_, new_n3725_})
2'b01 : new_n5211_ = 1'b1;
default : new_n5211_ = 1'b0;
endcase
casez ({new_n544_, new_n3726_})
2'b01 : new_n5212_ = 1'b1;
default : new_n5212_ = 1'b0;
endcase
casez ({new_n2922_, new_n3738_})
2'b01 : new_n5213_ = 1'b1;
default : new_n5213_ = 1'b0;
endcase
casez ({new_n193_, new_n279_, new_n1061_})
3'b11? : new_n5214_ = 1'b1;
3'b??1 : new_n5214_ = 1'b1;
default : new_n5214_ = 1'b0;
endcase
casez ({new_n1485_, new_n1716_})
2'b00 : new_n5215_ = 1'b1;
default : new_n5215_ = 1'b0;
endcase
casez ({new_n3519_, new_n3748_})
2'b01 : new_n5216_ = 1'b1;
default : new_n5216_ = 1'b0;
endcase
casez ({new_n657_, new_n3750_})
2'b01 : new_n5217_ = 1'b1;
default : new_n5217_ = 1'b0;
endcase
casez ({new_n949_, new_n1716_})
2'b00 : new_n5218_ = 1'b1;
default : new_n5218_ = 1'b0;
endcase
casez ({new_n91_, new_n680_, new_n1062_})
3'b11? : new_n5219_ = 1'b1;
3'b??1 : new_n5219_ = 1'b1;
default : new_n5219_ = 1'b0;
endcase
casez ({new_n1626_, new_n3755_})
2'b01 : new_n5220_ = 1'b1;
default : new_n5220_ = 1'b0;
endcase
casez ({new_n457_, new_n3764_})
2'b01 : new_n5221_ = 1'b1;
default : new_n5221_ = 1'b0;
endcase
casez ({new_n3085_, new_n3767_})
2'b01 : new_n5222_ = 1'b1;
default : new_n5222_ = 1'b0;
endcase
casez ({new_n2768_, new_n3773_})
2'b01 : new_n5223_ = 1'b1;
default : new_n5223_ = 1'b0;
endcase
casez ({new_n716_, new_n3775_})
2'b01 : new_n5224_ = 1'b1;
default : new_n5224_ = 1'b0;
endcase
casez ({new_n1070_, new_n1718_})
2'b00 : new_n5225_ = 1'b1;
default : new_n5225_ = 1'b0;
endcase
casez ({new_n1370_, new_n3779_})
2'b01 : new_n5226_ = 1'b1;
default : new_n5226_ = 1'b0;
endcase
casez ({new_n943_, new_n3783_})
2'b01 : new_n5227_ = 1'b1;
default : new_n5227_ = 1'b0;
endcase
casez ({new_n98_, new_n1064_, new_n329_, new_n654_})
4'b11?? : new_n5228_ = 1'b1;
4'b??11 : new_n5228_ = 1'b1;
default : new_n5228_ = 1'b0;
endcase
casez ({new_n724_, new_n1064_})
2'b00 : new_n5229_ = 1'b1;
default : new_n5229_ = 1'b0;
endcase
casez ({new_n1149_, new_n1723_})
2'b00 : new_n5230_ = 1'b1;
default : new_n5230_ = 1'b0;
endcase
casez ({new_n1464_, new_n1724_})
2'b00 : new_n5231_ = 1'b1;
default : new_n5231_ = 1'b0;
endcase
casez ({new_n908_, new_n1065_})
2'b00 : new_n5232_ = 1'b1;
default : new_n5232_ = 1'b0;
endcase
casez ({new_n613_, new_n3825_})
2'b01 : new_n5233_ = 1'b1;
default : new_n5233_ = 1'b0;
endcase
casez ({new_n1397_, new_n3827_})
2'b01 : new_n5234_ = 1'b1;
default : new_n5234_ = 1'b0;
endcase
casez ({u[1], new_n339_, new_n1066_})
3'b01? : new_n5235_ = 1'b1;
3'b??1 : new_n5235_ = 1'b1;
default : new_n5235_ = 1'b0;
endcase
casez ({new_n813_, new_n1728_})
2'b00 : new_n5236_ = 1'b1;
default : new_n5236_ = 1'b0;
endcase
casez ({new_n1209_, new_n1728_})
2'b00 : new_n5237_ = 1'b1;
default : new_n5237_ = 1'b0;
endcase
casez ({new_n2137_, new_n3842_})
2'b01 : new_n5238_ = 1'b1;
default : new_n5238_ = 1'b0;
endcase
casez ({new_n678_, new_n1067_})
2'b00 : new_n5239_ = 1'b1;
default : new_n5239_ = 1'b0;
endcase
casez ({new_n2156_, new_n3851_})
2'b01 : new_n5240_ = 1'b1;
default : new_n5240_ = 1'b0;
endcase
casez ({new_n2147_, new_n3855_})
2'b01 : new_n5241_ = 1'b1;
default : new_n5241_ = 1'b0;
endcase
casez ({new_n1593_, new_n3858_})
2'b01 : new_n5242_ = 1'b1;
default : new_n5242_ = 1'b0;
endcase
casez ({new_n830_, new_n1731_})
2'b00 : new_n5243_ = 1'b1;
default : new_n5243_ = 1'b0;
endcase
casez ({new_n1482_, new_n3864_})
2'b01 : new_n5244_ = 1'b1;
default : new_n5244_ = 1'b0;
endcase
casez ({new_n1061_, new_n1732_})
2'b00 : new_n5245_ = 1'b1;
default : new_n5245_ = 1'b0;
endcase
casez ({new_n1599_, new_n3867_})
2'b01 : new_n5246_ = 1'b1;
default : new_n5246_ = 1'b0;
endcase
casez ({new_n2808_, new_n3870_})
2'b01 : new_n5247_ = 1'b1;
default : new_n5247_ = 1'b0;
endcase
casez ({new_n1838_, new_n3875_})
2'b01 : new_n5248_ = 1'b1;
default : new_n5248_ = 1'b0;
endcase
casez ({new_n520_, new_n1069_})
2'b00 : new_n5249_ = 1'b1;
default : new_n5249_ = 1'b0;
endcase
casez ({new_n877_, new_n1733_})
2'b10 : new_n5250_ = 1'b1;
default : new_n5250_ = 1'b0;
endcase
casez ({new_n3499_, new_n3884_})
2'b01 : new_n5251_ = 1'b1;
default : new_n5251_ = 1'b0;
endcase
casez ({new_n977_, new_n1069_})
2'b00 : new_n5252_ = 1'b1;
default : new_n5252_ = 1'b0;
endcase
casez ({new_n96_, new_n345_, new_n3888_})
3'b01? : new_n5253_ = 1'b1;
3'b??0 : new_n5253_ = 1'b1;
default : new_n5253_ = 1'b0;
endcase
casez ({new_n520_, new_n3891_})
2'b01 : new_n5254_ = 1'b1;
default : new_n5254_ = 1'b0;
endcase
casez ({new_n237_, new_n783_, new_n1735_})
3'b11? : new_n5255_ = 1'b1;
3'b??1 : new_n5255_ = 1'b1;
default : new_n5255_ = 1'b0;
endcase
casez ({new_n901_, new_n3895_})
2'b01 : new_n5256_ = 1'b1;
default : new_n5256_ = 1'b0;
endcase
casez ({new_n419_, new_n3897_})
2'b01 : new_n5257_ = 1'b1;
default : new_n5257_ = 1'b0;
endcase
casez ({new_n1055_, new_n3902_})
2'b01 : new_n5258_ = 1'b1;
default : new_n5258_ = 1'b0;
endcase
casez ({new_n824_, new_n1737_})
2'b00 : new_n5259_ = 1'b1;
default : new_n5259_ = 1'b0;
endcase
casez ({new_n1585_, new_n1737_})
2'b00 : new_n5260_ = 1'b1;
default : new_n5260_ = 1'b0;
endcase
casez ({new_n1206_, new_n1738_})
2'b00 : new_n5261_ = 1'b1;
default : new_n5261_ = 1'b0;
endcase
casez ({new_n283_, new_n3920_})
2'b01 : new_n5262_ = 1'b1;
default : new_n5262_ = 1'b0;
endcase
casez ({new_n975_, new_n1740_})
2'b00 : new_n5263_ = 1'b1;
default : new_n5263_ = 1'b0;
endcase
casez ({new_n631_, new_n1740_})
2'b00 : new_n5264_ = 1'b1;
default : new_n5264_ = 1'b0;
endcase
casez ({new_n986_, new_n1740_})
2'b00 : new_n5265_ = 1'b1;
default : new_n5265_ = 1'b0;
endcase
casez ({new_n1634_, new_n3936_})
2'b01 : new_n5266_ = 1'b1;
default : new_n5266_ = 1'b0;
endcase
casez ({new_n1719_, new_n1741_})
2'b00 : new_n5267_ = 1'b1;
default : new_n5267_ = 1'b0;
endcase
casez ({new_n642_, new_n1072_})
2'b00 : new_n5268_ = 1'b1;
default : new_n5268_ = 1'b0;
endcase
casez ({new_n830_, new_n1742_})
2'b00 : new_n5269_ = 1'b1;
default : new_n5269_ = 1'b0;
endcase
casez ({new_n985_, new_n1742_})
2'b00 : new_n5270_ = 1'b1;
default : new_n5270_ = 1'b0;
endcase
casez ({new_n573_, new_n1742_})
2'b00 : new_n5271_ = 1'b1;
default : new_n5271_ = 1'b0;
endcase
casez ({new_n2148_, new_n3952_})
2'b01 : new_n5272_ = 1'b1;
default : new_n5272_ = 1'b0;
endcase
casez ({new_n83_, new_n629_, new_n3955_})
3'b10? : new_n5273_ = 1'b1;
3'b??0 : new_n5273_ = 1'b1;
default : new_n5273_ = 1'b0;
endcase
casez ({new_n3253_, new_n3961_})
2'b01 : new_n5274_ = 1'b1;
default : new_n5274_ = 1'b0;
endcase
casez ({new_n91_, new_n1744_, new_n146_, new_n294_})
4'b11?? : new_n5275_ = 1'b1;
4'b??11 : new_n5275_ = 1'b1;
default : new_n5275_ = 1'b0;
endcase
casez ({new_n3081_, new_n3964_})
2'b01 : new_n5276_ = 1'b1;
default : new_n5276_ = 1'b0;
endcase
casez ({x[0], new_n517_, new_n726_})
3'b01? : new_n5277_ = 1'b1;
3'b??1 : new_n5277_ = 1'b1;
default : new_n5277_ = 1'b0;
endcase
casez ({new_n2759_, new_n3967_})
2'b01 : new_n5278_ = 1'b1;
default : new_n5278_ = 1'b0;
endcase
casez ({new_n2101_, new_n3976_})
2'b11 : new_n5279_ = 1'b1;
default : new_n5279_ = 1'b0;
endcase
casez ({new_n1484_, new_n3977_})
2'b01 : new_n5280_ = 1'b1;
default : new_n5280_ = 1'b0;
endcase
casez ({new_n2640_, new_n3983_})
2'b01 : new_n5281_ = 1'b1;
default : new_n5281_ = 1'b0;
endcase
casez ({new_n988_, new_n1747_})
2'b00 : new_n5282_ = 1'b1;
default : new_n5282_ = 1'b0;
endcase
casez ({new_n402_, new_n3986_})
2'b01 : new_n5283_ = 1'b1;
default : new_n5283_ = 1'b0;
endcase
casez ({new_n1864_, new_n3989_})
2'b01 : new_n5284_ = 1'b1;
default : new_n5284_ = 1'b0;
endcase
casez ({new_n1208_, new_n1749_})
2'b00 : new_n5285_ = 1'b1;
default : new_n5285_ = 1'b0;
endcase
casez ({new_n482_, new_n1749_})
2'b00 : new_n5286_ = 1'b1;
default : new_n5286_ = 1'b0;
endcase
casez ({new_n3012_, new_n4000_})
2'b01 : new_n5287_ = 1'b1;
default : new_n5287_ = 1'b0;
endcase
casez ({new_n192_, new_n728_, new_n283_})
3'b11? : new_n5288_ = 1'b1;
3'b??1 : new_n5288_ = 1'b1;
default : new_n5288_ = 1'b0;
endcase
casez ({new_n974_, new_n4006_})
2'b01 : new_n5289_ = 1'b1;
default : new_n5289_ = 1'b0;
endcase
casez ({new_n720_, new_n4009_})
2'b11 : new_n5290_ = 1'b1;
default : new_n5290_ = 1'b0;
endcase
casez ({new_n3285_, new_n4011_})
2'b01 : new_n5291_ = 1'b1;
default : new_n5291_ = 1'b0;
endcase
casez ({new_n944_, new_n1751_})
2'b00 : new_n5292_ = 1'b1;
default : new_n5292_ = 1'b0;
endcase
casez ({new_n462_, new_n1752_})
2'b00 : new_n5293_ = 1'b1;
default : new_n5293_ = 1'b0;
endcase
casez ({new_n484_, new_n1752_})
2'b00 : new_n5294_ = 1'b1;
default : new_n5294_ = 1'b0;
endcase
casez ({new_n2634_, new_n4019_})
2'b01 : new_n5295_ = 1'b1;
default : new_n5295_ = 1'b0;
endcase
casez ({new_n722_, new_n1752_})
2'b00 : new_n5296_ = 1'b1;
default : new_n5296_ = 1'b0;
endcase
casez ({new_n727_, new_n4022_})
2'b01 : new_n5297_ = 1'b1;
default : new_n5297_ = 1'b0;
endcase
casez ({new_n1112_, new_n4029_})
2'b01 : new_n5298_ = 1'b1;
default : new_n5298_ = 1'b0;
endcase
casez ({new_n866_, new_n1753_})
2'b00 : new_n5299_ = 1'b1;
default : new_n5299_ = 1'b0;
endcase
casez ({new_n544_, new_n4030_})
2'b01 : new_n5300_ = 1'b1;
default : new_n5300_ = 1'b0;
endcase
casez ({new_n3470_, new_n4045_})
2'b01 : new_n5301_ = 1'b1;
default : new_n5301_ = 1'b0;
endcase
casez ({new_n2647_, new_n4049_})
2'b01 : new_n5302_ = 1'b1;
default : new_n5302_ = 1'b0;
endcase
casez ({new_n3368_, new_n4050_})
2'b01 : new_n5303_ = 1'b1;
default : new_n5303_ = 1'b0;
endcase
casez ({new_n1227_, new_n4059_})
2'b01 : new_n5304_ = 1'b1;
default : new_n5304_ = 1'b0;
endcase
casez ({new_n613_, new_n4070_})
2'b01 : new_n5305_ = 1'b1;
default : new_n5305_ = 1'b0;
endcase
casez ({new_n1480_, new_n4072_})
2'b01 : new_n5306_ = 1'b1;
default : new_n5306_ = 1'b0;
endcase
casez ({new_n4007_, new_n4074_})
2'b11 : new_n5307_ = 1'b1;
default : new_n5307_ = 1'b0;
endcase
casez ({new_n1218_, new_n4077_})
2'b01 : new_n5308_ = 1'b1;
default : new_n5308_ = 1'b0;
endcase
casez ({new_n1601_, new_n4085_})
2'b01 : new_n5309_ = 1'b1;
default : new_n5309_ = 1'b0;
endcase
casez ({new_n834_, new_n4088_})
2'b01 : new_n5310_ = 1'b1;
default : new_n5310_ = 1'b0;
endcase
casez ({new_n3514_, new_n4094_})
2'b01 : new_n5311_ = 1'b1;
default : new_n5311_ = 1'b0;
endcase
casez ({new_n97_, new_n297_, new_n4097_})
3'b11? : new_n5312_ = 1'b1;
3'b??0 : new_n5312_ = 1'b1;
default : new_n5312_ = 1'b0;
endcase
casez ({new_n4062_, new_n4106_})
2'b11 : new_n5313_ = 1'b1;
default : new_n5313_ = 1'b0;
endcase
casez ({new_n4005_, new_n4107_})
2'b11 : new_n5314_ = 1'b1;
default : new_n5314_ = 1'b0;
endcase
casez ({new_n1467_, new_n4108_})
2'b01 : new_n5315_ = 1'b1;
default : new_n5315_ = 1'b0;
endcase
casez ({new_n3107_, new_n4116_})
2'b01 : new_n5316_ = 1'b1;
default : new_n5316_ = 1'b0;
endcase
casez ({new_n645_, new_n4122_})
2'b01 : new_n5317_ = 1'b1;
default : new_n5317_ = 1'b0;
endcase
casez ({new_n3385_, new_n4124_})
2'b01 : new_n5318_ = 1'b1;
default : new_n5318_ = 1'b0;
endcase
casez ({new_n435_, new_n4126_})
2'b01 : new_n5319_ = 1'b1;
default : new_n5319_ = 1'b0;
endcase
casez ({new_n977_, new_n4128_})
2'b01 : new_n5320_ = 1'b1;
default : new_n5320_ = 1'b0;
endcase
casez ({new_n1734_, new_n4132_})
2'b01 : new_n5321_ = 1'b1;
default : new_n5321_ = 1'b0;
endcase
casez ({new_n3511_, new_n4134_})
2'b01 : new_n5322_ = 1'b1;
default : new_n5322_ = 1'b0;
endcase
casez ({new_n816_, new_n4138_})
2'b01 : new_n5323_ = 1'b1;
default : new_n5323_ = 1'b0;
endcase
casez ({new_n2832_, new_n4151_})
2'b01 : new_n5324_ = 1'b1;
default : new_n5324_ = 1'b0;
endcase
casez ({new_n429_, new_n4163_})
2'b01 : new_n5325_ = 1'b1;
default : new_n5325_ = 1'b0;
endcase
casez ({new_n4113_, new_n4166_})
2'b11 : new_n5326_ = 1'b1;
default : new_n5326_ = 1'b0;
endcase
casez ({new_n94_, new_n98_, new_n4178_})
3'b11? : new_n5327_ = 1'b1;
3'b??0 : new_n5327_ = 1'b1;
default : new_n5327_ = 1'b0;
endcase
casez ({new_n3333_, new_n4180_})
2'b01 : new_n5328_ = 1'b1;
default : new_n5328_ = 1'b0;
endcase
casez ({new_n322_, new_n4181_})
2'b01 : new_n5329_ = 1'b1;
default : new_n5329_ = 1'b0;
endcase
casez ({new_n2154_, new_n4187_})
2'b01 : new_n5330_ = 1'b1;
default : new_n5330_ = 1'b0;
endcase
casez ({new_n4052_, new_n4189_})
2'b11 : new_n5331_ = 1'b1;
default : new_n5331_ = 1'b0;
endcase
casez ({new_n1831_, new_n4190_})
2'b01 : new_n5332_ = 1'b1;
default : new_n5332_ = 1'b0;
endcase
casez ({new_n170_, new_n2786_, new_n4216_})
3'b10? : new_n5333_ = 1'b1;
3'b??0 : new_n5333_ = 1'b1;
default : new_n5333_ = 1'b0;
endcase
casez ({new_n1070_, new_n1105_})
2'b00 : new_n5334_ = 1'b1;
default : new_n5334_ = 1'b0;
endcase
casez ({new_n3716_, new_n4225_})
2'b11 : new_n5335_ = 1'b1;
default : new_n5335_ = 1'b0;
endcase
casez ({new_n270_, new_n4227_})
2'b01 : new_n5336_ = 1'b1;
default : new_n5336_ = 1'b0;
endcase
casez ({new_n840_, new_n4232_})
2'b01 : new_n5337_ = 1'b1;
default : new_n5337_ = 1'b0;
endcase
casez ({new_n3134_, new_n4238_})
2'b01 : new_n5338_ = 1'b1;
default : new_n5338_ = 1'b0;
endcase
casez ({new_n3538_, new_n4239_})
2'b01 : new_n5339_ = 1'b1;
default : new_n5339_ = 1'b0;
endcase
casez ({new_n1631_, new_n4243_})
2'b01 : new_n5340_ = 1'b1;
default : new_n5340_ = 1'b0;
endcase
casez ({new_n838_, new_n4246_})
2'b01 : new_n5341_ = 1'b1;
default : new_n5341_ = 1'b0;
endcase
casez ({new_n246_, new_n388_, new_n4250_})
3'b11? : new_n5342_ = 1'b1;
3'b??0 : new_n5342_ = 1'b1;
default : new_n5342_ = 1'b0;
endcase
casez ({new_n1327_, new_n4257_})
2'b01 : new_n5343_ = 1'b1;
default : new_n5343_ = 1'b0;
endcase
casez ({new_n1616_, new_n4272_})
2'b01 : new_n5344_ = 1'b1;
default : new_n5344_ = 1'b0;
endcase
casez ({new_n79_, new_n2784_, new_n4278_})
3'b10? : new_n5345_ = 1'b1;
3'b??0 : new_n5345_ = 1'b1;
default : new_n5345_ = 1'b0;
endcase
casez ({new_n808_, new_n4286_})
2'b01 : new_n5346_ = 1'b1;
default : new_n5346_ = 1'b0;
endcase
casez ({new_n1111_, new_n4295_})
2'b01 : new_n5347_ = 1'b1;
default : new_n5347_ = 1'b0;
endcase
casez ({new_n3204_, new_n4296_})
2'b01 : new_n5348_ = 1'b1;
default : new_n5348_ = 1'b0;
endcase
casez ({new_n1225_, new_n4297_})
2'b01 : new_n5349_ = 1'b1;
default : new_n5349_ = 1'b0;
endcase
casez ({new_n3343_, new_n4299_})
2'b01 : new_n5350_ = 1'b1;
default : new_n5350_ = 1'b0;
endcase
casez ({new_n1136_, new_n4300_})
2'b01 : new_n5351_ = 1'b1;
default : new_n5351_ = 1'b0;
endcase
casez ({new_n1479_, new_n4302_})
2'b01 : new_n5352_ = 1'b1;
default : new_n5352_ = 1'b0;
endcase
casez ({new_n699_, new_n4321_})
2'b01 : new_n5353_ = 1'b1;
default : new_n5353_ = 1'b0;
endcase
casez ({new_n3175_, new_n4327_})
2'b01 : new_n5354_ = 1'b1;
default : new_n5354_ = 1'b0;
endcase
casez ({new_n1631_, new_n4332_})
2'b01 : new_n5355_ = 1'b1;
default : new_n5355_ = 1'b0;
endcase
casez ({new_n1203_, new_n1823_})
2'b00 : new_n5356_ = 1'b1;
default : new_n5356_ = 1'b0;
endcase
casez ({new_n2144_, new_n4339_})
2'b01 : new_n5357_ = 1'b1;
default : new_n5357_ = 1'b0;
endcase
casez ({new_n831_, new_n4342_})
2'b01 : new_n5358_ = 1'b1;
default : new_n5358_ = 1'b0;
endcase
casez ({new_n2069_, new_n4346_})
2'b11 : new_n5359_ = 1'b1;
default : new_n5359_ = 1'b0;
endcase
casez ({new_n1325_, new_n4352_})
2'b01 : new_n5360_ = 1'b1;
default : new_n5360_ = 1'b0;
endcase
casez ({new_n402_, new_n4354_})
2'b01 : new_n5361_ = 1'b1;
default : new_n5361_ = 1'b0;
endcase
casez ({new_n3154_, new_n4356_})
2'b01 : new_n5362_ = 1'b1;
default : new_n5362_ = 1'b0;
endcase
casez ({new_n2791_, new_n4363_})
2'b01 : new_n5363_ = 1'b1;
default : new_n5363_ = 1'b0;
endcase
casez ({new_n3027_, new_n4365_})
2'b01 : new_n5364_ = 1'b1;
default : new_n5364_ = 1'b0;
endcase
casez ({new_n573_, new_n4368_})
2'b01 : new_n5365_ = 1'b1;
default : new_n5365_ = 1'b0;
endcase
casez ({new_n1751_, new_n1829_})
2'b00 : new_n5366_ = 1'b1;
default : new_n5366_ = 1'b0;
endcase
casez ({new_n756_, new_n4371_})
2'b01 : new_n5367_ = 1'b1;
default : new_n5367_ = 1'b0;
endcase
casez ({new_n1826_, new_n4372_})
2'b01 : new_n5368_ = 1'b1;
default : new_n5368_ = 1'b0;
endcase
casez ({new_n1274_, new_n4375_})
2'b01 : new_n5369_ = 1'b1;
default : new_n5369_ = 1'b0;
endcase
casez ({new_n726_, new_n4378_})
2'b01 : new_n5370_ = 1'b1;
default : new_n5370_ = 1'b0;
endcase
casez ({new_n1220_, new_n1830_})
2'b00 : new_n5371_ = 1'b1;
default : new_n5371_ = 1'b0;
endcase
casez ({new_n720_, new_n1115_})
2'b10 : new_n5372_ = 1'b1;
default : new_n5372_ = 1'b0;
endcase
casez ({new_n973_, new_n1832_})
2'b00 : new_n5373_ = 1'b1;
default : new_n5373_ = 1'b0;
endcase
casez ({new_n3153_, new_n4391_})
2'b01 : new_n5374_ = 1'b1;
default : new_n5374_ = 1'b0;
endcase
casez ({new_n1042_, new_n4392_})
2'b01 : new_n5375_ = 1'b1;
default : new_n5375_ = 1'b0;
endcase
casez ({new_n755_, new_n1832_})
2'b00 : new_n5376_ = 1'b1;
default : new_n5376_ = 1'b0;
endcase
casez ({new_n376_, new_n462_})
2'b00 : new_n5377_ = 1'b1;
default : new_n5377_ = 1'b0;
endcase
casez ({new_n1722_, new_n4403_})
2'b01 : new_n5378_ = 1'b1;
default : new_n5378_ = 1'b0;
endcase
casez ({new_n988_, new_n4411_})
2'b01 : new_n5379_ = 1'b1;
default : new_n5379_ = 1'b0;
endcase
casez ({new_n624_, new_n4422_})
2'b01 : new_n5380_ = 1'b1;
default : new_n5380_ = 1'b0;
endcase
casez ({new_n3694_, new_n4430_})
2'b11 : new_n5381_ = 1'b1;
default : new_n5381_ = 1'b0;
endcase
casez ({new_n1497_, new_n4436_})
2'b01 : new_n5382_ = 1'b1;
default : new_n5382_ = 1'b0;
endcase
casez ({new_n4426_, new_n4441_})
2'b11 : new_n5383_ = 1'b1;
default : new_n5383_ = 1'b0;
endcase
casez ({new_n756_, new_n1839_})
2'b00 : new_n5384_ = 1'b1;
default : new_n5384_ = 1'b0;
endcase
casez ({new_n727_, new_n4448_})
2'b01 : new_n5385_ = 1'b1;
default : new_n5385_ = 1'b0;
endcase
casez ({new_n727_, new_n1842_})
2'b00 : new_n5386_ = 1'b1;
default : new_n5386_ = 1'b0;
endcase
casez ({new_n582_, new_n4467_})
2'b01 : new_n5387_ = 1'b1;
default : new_n5387_ = 1'b0;
endcase
casez ({new_n464_, new_n1845_})
2'b00 : new_n5388_ = 1'b1;
default : new_n5388_ = 1'b0;
endcase
casez ({new_n477_, new_n1846_})
2'b00 : new_n5389_ = 1'b1;
default : new_n5389_ = 1'b0;
endcase
casez ({new_n903_, new_n4488_})
2'b01 : new_n5390_ = 1'b1;
default : new_n5390_ = 1'b0;
endcase
casez ({new_n3165_, new_n4490_})
2'b01 : new_n5391_ = 1'b1;
default : new_n5391_ = 1'b0;
endcase
casez ({new_n1482_, new_n4502_})
2'b01 : new_n5392_ = 1'b1;
default : new_n5392_ = 1'b0;
endcase
casez ({new_n568_, new_n1122_})
2'b00 : new_n5393_ = 1'b1;
default : new_n5393_ = 1'b0;
endcase
casez ({new_n903_, new_n4503_})
2'b01 : new_n5394_ = 1'b1;
default : new_n5394_ = 1'b0;
endcase
casez ({new_n263_, new_n321_, new_n750_})
3'b11? : new_n5395_ = 1'b1;
3'b??1 : new_n5395_ = 1'b1;
default : new_n5395_ = 1'b0;
endcase
casez ({new_n98_, new_n1850_, new_n646_})
3'b11? : new_n5396_ = 1'b1;
3'b??1 : new_n5396_ = 1'b1;
default : new_n5396_ = 1'b0;
endcase
casez ({new_n1755_, new_n4519_})
2'b01 : new_n5397_ = 1'b1;
default : new_n5397_ = 1'b0;
endcase
casez ({new_n3000_, new_n4526_})
2'b01 : new_n5398_ = 1'b1;
default : new_n5398_ = 1'b0;
endcase
casez ({new_n1749_, new_n1853_})
2'b00 : new_n5399_ = 1'b1;
default : new_n5399_ = 1'b0;
endcase
casez ({new_n426_, new_n751_})
2'b00 : new_n5400_ = 1'b1;
default : new_n5400_ = 1'b0;
endcase
casez ({new_n2148_, new_n4533_})
2'b01 : new_n5401_ = 1'b1;
default : new_n5401_ = 1'b0;
endcase
casez ({new_n906_, new_n4535_})
2'b01 : new_n5402_ = 1'b1;
default : new_n5402_ = 1'b0;
endcase
casez ({new_n92_, new_n467_, new_n93_, new_n312_})
4'b11?? : new_n5403_ = 1'b1;
4'b??11 : new_n5403_ = 1'b1;
default : new_n5403_ = 1'b0;
endcase
casez ({new_n2116_, new_n4537_})
2'b01 : new_n5404_ = 1'b1;
default : new_n5404_ = 1'b0;
endcase
casez ({new_n2160_, new_n4541_})
2'b01 : new_n5405_ = 1'b1;
default : new_n5405_ = 1'b0;
endcase
casez ({new_n1492_, new_n4543_})
2'b01 : new_n5406_ = 1'b1;
default : new_n5406_ = 1'b0;
endcase
casez ({new_n426_, new_n1125_})
2'b00 : new_n5407_ = 1'b1;
default : new_n5407_ = 1'b0;
endcase
casez ({new_n1460_, new_n4548_})
2'b01 : new_n5408_ = 1'b1;
default : new_n5408_ = 1'b0;
endcase
casez ({new_n905_, new_n4549_})
2'b01 : new_n5409_ = 1'b1;
default : new_n5409_ = 1'b0;
endcase
casez ({new_n665_, new_n1857_})
2'b00 : new_n5410_ = 1'b1;
default : new_n5410_ = 1'b0;
endcase
casez ({new_n756_, new_n4561_})
2'b01 : new_n5411_ = 1'b1;
default : new_n5411_ = 1'b0;
endcase
casez ({new_n1478_, new_n1857_})
2'b00 : new_n5412_ = 1'b1;
default : new_n5412_ = 1'b0;
endcase
casez ({new_n664_, new_n4564_})
2'b01 : new_n5413_ = 1'b1;
default : new_n5413_ = 1'b0;
endcase
casez ({new_n3220_, new_n4565_})
2'b01 : new_n5414_ = 1'b1;
default : new_n5414_ = 1'b0;
endcase
casez ({new_n1314_, new_n4567_})
2'b01 : new_n5415_ = 1'b1;
default : new_n5415_ = 1'b0;
endcase
casez ({new_n1056_, new_n4568_})
2'b01 : new_n5416_ = 1'b1;
default : new_n5416_ = 1'b0;
endcase
casez ({new_n976_, new_n4580_})
2'b00 : new_n5417_ = 1'b1;
default : new_n5417_ = 1'b0;
endcase
casez ({new_n1056_, new_n4592_})
2'b00 : new_n5418_ = 1'b1;
default : new_n5418_ = 1'b0;
endcase
casez ({new_n1215_, new_n1865_})
2'b00 : new_n5419_ = 1'b1;
default : new_n5419_ = 1'b0;
endcase
casez ({new_n2787_, new_n4619_})
2'b00 : new_n5420_ = 1'b1;
default : new_n5420_ = 1'b0;
endcase
casez ({new_n1470_, new_n4626_})
2'b00 : new_n5421_ = 1'b1;
default : new_n5421_ = 1'b0;
endcase
casez ({new_n1490_, new_n4629_})
2'b00 : new_n5422_ = 1'b1;
default : new_n5422_ = 1'b0;
endcase
casez ({new_n104_, new_n1872_, new_n1062_})
3'b11? : new_n5423_ = 1'b1;
3'b??1 : new_n5423_ = 1'b1;
default : new_n5423_ = 1'b0;
endcase
casez ({new_n997_, new_n1133_})
2'b00 : new_n5424_ = 1'b1;
default : new_n5424_ = 1'b0;
endcase
casez ({new_n1465_, new_n1877_})
2'b00 : new_n5425_ = 1'b1;
default : new_n5425_ = 1'b0;
endcase
casez ({new_n708_, new_n1137_})
2'b00 : new_n5426_ = 1'b1;
default : new_n5426_ = 1'b0;
endcase
casez ({y[2], new_n721_, new_n1138_})
3'b10? : new_n5427_ = 1'b1;
3'b??1 : new_n5427_ = 1'b1;
default : new_n5427_ = 1'b0;
endcase
casez ({new_n1215_, new_n1896_})
2'b00 : new_n5428_ = 1'b1;
default : new_n5428_ = 1'b0;
endcase
casez ({new_n905_, new_n1142_})
2'b00 : new_n5429_ = 1'b1;
default : new_n5429_ = 1'b0;
endcase
casez ({new_n245_, new_n479_})
2'b00 : new_n5430_ = 1'b1;
default : new_n5430_ = 1'b0;
endcase
casez ({new_n391_, new_n801_})
2'b10 : new_n5431_ = 1'b1;
default : new_n5431_ = 1'b0;
endcase
casez ({new_n385_, new_n1208_})
2'b11 : new_n5432_ = 1'b1;
default : new_n5432_ = 1'b0;
endcase
casez ({new_n223_, new_n1226_})
2'b11 : new_n5433_ = 1'b1;
default : new_n5433_ = 1'b0;
endcase
casez ({new_n96_, new_n2149_})
2'b11 : new_n5434_ = 1'b1;
default : new_n5434_ = 1'b0;
endcase
casez ({new_n97_, new_n2150_})
2'b11 : new_n5435_ = 1'b1;
default : new_n5435_ = 1'b0;
endcase
casez ({new_n257_, new_n846_})
2'b11 : new_n5436_ = 1'b1;
default : new_n5436_ = 1'b0;
endcase
casez ({new_n226_, new_n566_})
2'b11 : new_n5437_ = 1'b1;
default : new_n5437_ = 1'b0;
endcase
casez ({new_n151_, new_n610_})
2'b11 : new_n5438_ = 1'b1;
default : new_n5438_ = 1'b0;
endcase
casez ({new_n531_, new_n1470_})
2'b11 : new_n5439_ = 1'b1;
default : new_n5439_ = 1'b0;
endcase
casez ({new_n180_, new_n2805_})
2'b11 : new_n5440_ = 1'b1;
default : new_n5440_ = 1'b0;
endcase
casez ({new_n168_, new_n973_})
2'b11 : new_n5441_ = 1'b1;
default : new_n5441_ = 1'b0;
endcase
casez ({new_n139_, new_n2834_})
2'b11 : new_n5442_ = 1'b1;
default : new_n5442_ = 1'b0;
endcase
casez ({new_n459_, new_n982_})
2'b11 : new_n5443_ = 1'b1;
default : new_n5443_ = 1'b0;
endcase
casez ({new_n429_, new_n987_})
2'b11 : new_n5444_ = 1'b1;
default : new_n5444_ = 1'b0;
endcase
casez ({new_n423_, new_n987_})
2'b11 : new_n5445_ = 1'b1;
default : new_n5445_ = 1'b0;
endcase
casez ({new_n199_, new_n368_})
2'b11 : new_n5446_ = 1'b1;
default : new_n5446_ = 1'b0;
endcase
casez ({new_n270_, new_n675_})
2'b11 : new_n5447_ = 1'b1;
default : new_n5447_ = 1'b0;
endcase
casez ({new_n401_, new_n1060_})
2'b11 : new_n5448_ = 1'b1;
default : new_n5448_ = 1'b0;
endcase
casez ({new_n358_, new_n1746_})
2'b11 : new_n5449_ = 1'b1;
default : new_n5449_ = 1'b0;
endcase
casez ({new_n234_, new_n733_})
2'b11 : new_n5450_ = 1'b1;
default : new_n5450_ = 1'b0;
endcase
casez ({new_n757_, new_n1797_})
2'b11 : new_n5451_ = 1'b1;
default : new_n5451_ = 1'b0;
endcase
casez ({new_n159_, new_n754_})
2'b11 : new_n5452_ = 1'b1;
default : new_n5452_ = 1'b0;
endcase
casez ({new_n93_, new_n270_})
2'b11 : new_n5453_ = 1'b1;
default : new_n5453_ = 1'b0;
endcase
casez ({new_n285_, new_n561_})
2'b11 : new_n5454_ = 1'b1;
default : new_n5454_ = 1'b0;
endcase
casez ({new_n207_, new_n611_})
2'b11 : new_n5455_ = 1'b1;
default : new_n5455_ = 1'b0;
endcase
casez ({new_n182_, new_n625_})
2'b11 : new_n5456_ = 1'b1;
default : new_n5456_ = 1'b0;
endcase
casez ({new_n134_, new_n463_})
2'b11 : new_n5457_ = 1'b1;
default : new_n5457_ = 1'b0;
endcase
casez ({new_n115_, new_n246_})
2'b11 : new_n5458_ = 1'b1;
default : new_n5458_ = 1'b0;
endcase
casez ({new_n819_, new_n1143_})
2'b00 : new_n5459_ = 1'b1;
default : new_n5459_ = 1'b0;
endcase
casez ({new_n1452_, new_n1915_})
2'b00 : new_n5460_ = 1'b1;
default : new_n5460_ = 1'b0;
endcase
casez ({new_n4377_, new_n4857_})
2'b11 : new_n5461_ = 1'b1;
default : new_n5461_ = 1'b0;
endcase
casez ({new_n697_, new_n4860_})
2'b01 : new_n5462_ = 1'b1;
default : new_n5462_ = 1'b0;
endcase
casez ({new_n2802_, new_n4861_})
2'b01 : new_n5463_ = 1'b1;
default : new_n5463_ = 1'b0;
endcase
casez ({new_n4221_, new_n4862_})
2'b11 : new_n5464_ = 1'b1;
default : new_n5464_ = 1'b0;
endcase
casez ({new_n84_, new_n277_, new_n4863_})
3'b01? : new_n5465_ = 1'b1;
3'b??0 : new_n5465_ = 1'b1;
default : new_n5465_ = 1'b0;
endcase
casez ({new_n1028_, new_n4864_})
2'b01 : new_n5466_ = 1'b1;
default : new_n5466_ = 1'b0;
endcase
casez ({new_n365_, new_n4884_})
2'b01 : new_n5467_ = 1'b1;
default : new_n5467_ = 1'b0;
endcase
casez ({new_n3840_, new_n4886_})
2'b01 : new_n5468_ = 1'b1;
default : new_n5468_ = 1'b0;
endcase
casez ({new_n3019_, new_n4892_})
2'b01 : new_n5469_ = 1'b1;
default : new_n5469_ = 1'b0;
endcase
casez ({new_n547_, new_n4899_})
2'b01 : new_n5470_ = 1'b1;
default : new_n5470_ = 1'b0;
endcase
casez ({new_n4036_, new_n4906_})
2'b11 : new_n5471_ = 1'b1;
default : new_n5471_ = 1'b0;
endcase
casez ({new_n3972_, new_n4909_})
2'b11 : new_n5472_ = 1'b1;
default : new_n5472_ = 1'b0;
endcase
casez ({new_n546_, new_n4916_})
2'b01 : new_n5473_ = 1'b1;
default : new_n5473_ = 1'b0;
endcase
casez ({new_n84_, new_n1775_, new_n4918_})
3'b10? : new_n5474_ = 1'b1;
3'b??0 : new_n5474_ = 1'b1;
default : new_n5474_ = 1'b0;
endcase
casez ({new_n3647_, new_n4919_})
2'b01 : new_n5475_ = 1'b1;
default : new_n5475_ = 1'b0;
endcase
casez ({new_n1487_, new_n4927_})
2'b01 : new_n5476_ = 1'b1;
default : new_n5476_ = 1'b0;
endcase
casez ({new_n4172_, new_n4929_})
2'b11 : new_n5477_ = 1'b1;
default : new_n5477_ = 1'b0;
endcase
casez ({new_n3865_, new_n4930_})
2'b01 : new_n5478_ = 1'b1;
default : new_n5478_ = 1'b0;
endcase
casez ({new_n1755_, new_n4934_})
2'b01 : new_n5479_ = 1'b1;
default : new_n5479_ = 1'b0;
endcase
casez ({new_n2826_, new_n4935_})
2'b01 : new_n5480_ = 1'b1;
default : new_n5480_ = 1'b0;
endcase
casez ({new_n1559_, new_n4939_})
2'b01 : new_n5481_ = 1'b1;
default : new_n5481_ = 1'b0;
endcase
casez ({new_n4805_, new_n4942_})
2'b11 : new_n5482_ = 1'b1;
default : new_n5482_ = 1'b0;
endcase
casez ({new_n3868_, new_n4943_})
2'b01 : new_n5483_ = 1'b1;
default : new_n5483_ = 1'b0;
endcase
casez ({new_n2818_, new_n4955_})
2'b01 : new_n5484_ = 1'b1;
default : new_n5484_ = 1'b0;
endcase
casez ({new_n1847_, new_n4961_})
2'b01 : new_n5485_ = 1'b1;
default : new_n5485_ = 1'b0;
endcase
casez ({new_n4714_, new_n4962_})
2'b11 : new_n5486_ = 1'b1;
default : new_n5486_ = 1'b0;
endcase
casez ({new_n3953_, new_n4970_})
2'b01 : new_n5487_ = 1'b1;
default : new_n5487_ = 1'b0;
endcase
casez ({new_n2816_, new_n4971_})
2'b01 : new_n5488_ = 1'b1;
default : new_n5488_ = 1'b0;
endcase
casez ({new_n2816_, new_n4974_})
2'b01 : new_n5489_ = 1'b1;
default : new_n5489_ = 1'b0;
endcase
casez ({new_n2188_, new_n4990_})
2'b11 : new_n5490_ = 1'b1;
default : new_n5490_ = 1'b0;
endcase
casez ({new_n4033_, new_n4991_})
2'b01 : new_n5491_ = 1'b1;
default : new_n5491_ = 1'b0;
endcase
casez ({new_n670_, new_n4995_})
2'b01 : new_n5492_ = 1'b1;
default : new_n5492_ = 1'b0;
endcase
casez ({new_n1525_, new_n1928_})
2'b00 : new_n5493_ = 1'b1;
default : new_n5493_ = 1'b0;
endcase
casez ({new_n644_, new_n4998_})
2'b01 : new_n5494_ = 1'b1;
default : new_n5494_ = 1'b0;
endcase
casez ({new_n2831_, new_n5001_})
2'b01 : new_n5495_ = 1'b1;
default : new_n5495_ = 1'b0;
endcase
casez ({new_n5930_, new_n5004_})
2'b1? : new_n5496_ = 1'b1;
2'b?0 : new_n5496_ = 1'b1;
default : new_n5496_ = 1'b0;
endcase
casez ({new_n1738_, new_n5007_})
2'b01 : new_n5497_ = 1'b1;
default : new_n5497_ = 1'b0;
endcase
casez ({new_n1736_, new_n5011_})
2'b01 : new_n5498_ = 1'b1;
default : new_n5498_ = 1'b0;
endcase
casez ({new_n684_, new_n5014_})
2'b01 : new_n5499_ = 1'b1;
default : new_n5499_ = 1'b0;
endcase
casez ({new_n1674_, new_n5017_})
2'b01 : new_n5500_ = 1'b1;
default : new_n5500_ = 1'b0;
endcase
casez ({new_n2984_, new_n5019_})
2'b01 : new_n5501_ = 1'b1;
default : new_n5501_ = 1'b0;
endcase
casez ({new_n3549_, new_n5020_})
2'b01 : new_n5502_ = 1'b1;
default : new_n5502_ = 1'b0;
endcase
casez ({new_n1838_, new_n5040_})
2'b01 : new_n5503_ = 1'b1;
default : new_n5503_ = 1'b0;
endcase
casez ({new_n4084_, new_n5048_})
2'b11 : new_n5504_ = 1'b1;
default : new_n5504_ = 1'b0;
endcase
casez ({new_n3057_, new_n5049_})
2'b01 : new_n5505_ = 1'b1;
default : new_n5505_ = 1'b0;
endcase
casez ({new_n4027_, new_n5064_})
2'b11 : new_n5506_ = 1'b1;
default : new_n5506_ = 1'b0;
endcase
casez ({new_n2241_, new_n5066_})
2'b11 : new_n5507_ = 1'b1;
default : new_n5507_ = 1'b0;
endcase
casez ({new_n684_, new_n1934_})
2'b00 : new_n5508_ = 1'b1;
default : new_n5508_ = 1'b0;
endcase
casez ({new_n1473_, new_n5076_})
2'b01 : new_n5509_ = 1'b1;
default : new_n5509_ = 1'b0;
endcase
casez ({new_n841_, new_n5079_})
2'b01 : new_n5510_ = 1'b1;
default : new_n5510_ = 1'b0;
endcase
casez ({new_n3893_, new_n5085_})
2'b11 : new_n5511_ = 1'b1;
default : new_n5511_ = 1'b0;
endcase
casez ({new_n1712_, new_n5086_})
2'b01 : new_n5512_ = 1'b1;
default : new_n5512_ = 1'b0;
endcase
casez ({new_n4500_, new_n5088_})
2'b11 : new_n5513_ = 1'b1;
default : new_n5513_ = 1'b0;
endcase
casez ({new_n1414_, new_n5090_})
2'b01 : new_n5514_ = 1'b1;
default : new_n5514_ = 1'b0;
endcase
casez ({new_n164_, new_n728_, new_n5094_})
3'b11? : new_n5515_ = 1'b1;
3'b??0 : new_n5515_ = 1'b1;
default : new_n5515_ = 1'b0;
endcase
casez ({new_n4073_, new_n5104_})
2'b11 : new_n5516_ = 1'b1;
default : new_n5516_ = 1'b0;
endcase
casez ({new_n4241_, new_n5110_})
2'b11 : new_n5517_ = 1'b1;
default : new_n5517_ = 1'b0;
endcase
casez ({new_n1719_, new_n5113_})
2'b01 : new_n5518_ = 1'b1;
default : new_n5518_ = 1'b0;
endcase
casez ({new_n3945_, new_n5114_})
2'b01 : new_n5519_ = 1'b1;
default : new_n5519_ = 1'b0;
endcase
casez ({new_n3957_, new_n5115_})
2'b11 : new_n5520_ = 1'b1;
default : new_n5520_ = 1'b0;
endcase
casez ({new_n562_, new_n5118_})
2'b01 : new_n5521_ = 1'b1;
default : new_n5521_ = 1'b0;
endcase
casez ({new_n1686_, new_n5119_})
2'b01 : new_n5522_ = 1'b1;
default : new_n5522_ = 1'b0;
endcase
casez ({new_n1501_, new_n5129_})
2'b01 : new_n5523_ = 1'b1;
default : new_n5523_ = 1'b0;
endcase
casez ({new_n3803_, new_n5132_})
2'b01 : new_n5524_ = 1'b1;
default : new_n5524_ = 1'b0;
endcase
casez ({new_n1524_, new_n5133_})
2'b01 : new_n5525_ = 1'b1;
default : new_n5525_ = 1'b0;
endcase
casez ({new_n2194_, new_n5140_})
2'b11 : new_n5526_ = 1'b1;
default : new_n5526_ = 1'b0;
endcase
casez ({new_n4123_, new_n5142_})
2'b11 : new_n5527_ = 1'b1;
default : new_n5527_ = 1'b0;
endcase
casez ({new_n590_, new_n1164_})
2'b00 : new_n5528_ = 1'b1;
default : new_n5528_ = 1'b0;
endcase
casez ({new_n563_, new_n1165_})
2'b00 : new_n5529_ = 1'b1;
default : new_n5529_ = 1'b0;
endcase
casez ({new_n4171_, new_n5146_})
2'b01 : new_n5530_ = 1'b1;
default : new_n5530_ = 1'b0;
endcase
casez ({new_n4115_, new_n5147_})
2'b11 : new_n5531_ = 1'b1;
default : new_n5531_ = 1'b0;
endcase
casez ({new_n4722_, new_n5148_})
2'b11 : new_n5532_ = 1'b1;
default : new_n5532_ = 1'b0;
endcase
casez ({new_n4307_, new_n5153_})
2'b11 : new_n5533_ = 1'b1;
default : new_n5533_ = 1'b0;
endcase
casez ({new_n4341_, new_n5175_})
2'b11 : new_n5534_ = 1'b1;
default : new_n5534_ = 1'b0;
endcase
casez ({new_n916_, new_n5189_})
2'b01 : new_n5535_ = 1'b1;
default : new_n5535_ = 1'b0;
endcase
casez ({new_n1718_, new_n5191_})
2'b01 : new_n5536_ = 1'b1;
default : new_n5536_ = 1'b0;
endcase
casez ({new_n3892_, new_n5197_})
2'b01 : new_n5537_ = 1'b1;
default : new_n5537_ = 1'b0;
endcase
casez ({new_n4607_, new_n5199_})
2'b01 : new_n5538_ = 1'b1;
default : new_n5538_ = 1'b0;
endcase
casez ({new_n1666_, new_n5202_})
2'b01 : new_n5539_ = 1'b1;
default : new_n5539_ = 1'b0;
endcase
casez ({new_n917_, new_n5212_})
2'b01 : new_n5540_ = 1'b1;
default : new_n5540_ = 1'b0;
endcase
casez ({new_n1743_, new_n5217_})
2'b01 : new_n5541_ = 1'b1;
default : new_n5541_ = 1'b0;
endcase
casez ({new_n4625_, new_n5231_})
2'b01 : new_n5542_ = 1'b1;
default : new_n5542_ = 1'b0;
endcase
casez ({new_n4317_, new_n5238_})
2'b11 : new_n5543_ = 1'b1;
default : new_n5543_ = 1'b0;
endcase
casez ({new_n3915_, new_n5247_})
2'b01 : new_n5544_ = 1'b1;
default : new_n5544_ = 1'b0;
endcase
casez ({new_n3619_, new_n5254_})
2'b01 : new_n5545_ = 1'b1;
default : new_n5545_ = 1'b0;
endcase
casez ({new_n670_, new_n5261_})
2'b01 : new_n5546_ = 1'b1;
default : new_n5546_ = 1'b0;
endcase
casez ({new_n2336_, new_n5271_})
2'b01 : new_n5547_ = 1'b1;
default : new_n5547_ = 1'b0;
endcase
casez ({new_n4425_, new_n5283_})
2'b11 : new_n5548_ = 1'b1;
default : new_n5548_ = 1'b0;
endcase
casez ({new_n704_, new_n787_})
2'b00 : new_n5549_ = 1'b1;
default : new_n5549_ = 1'b0;
endcase
casez ({new_n410_, new_n1169_})
2'b10 : new_n5550_ = 1'b1;
default : new_n5550_ = 1'b0;
endcase
casez ({new_n5054_, new_n5300_})
2'b11 : new_n5551_ = 1'b1;
default : new_n5551_ = 1'b0;
endcase
casez ({new_n2282_, new_n5302_})
2'b11 : new_n5552_ = 1'b1;
default : new_n5552_ = 1'b0;
endcase
casez ({new_n1701_, new_n5306_})
2'b01 : new_n5553_ = 1'b1;
default : new_n5553_ = 1'b0;
endcase
casez ({new_n4081_, new_n5308_})
2'b11 : new_n5554_ = 1'b1;
default : new_n5554_ = 1'b0;
endcase
casez ({new_n546_, new_n5310_})
2'b01 : new_n5555_ = 1'b1;
default : new_n5555_ = 1'b0;
endcase
casez ({new_n5039_, new_n5314_})
2'b11 : new_n5556_ = 1'b1;
default : new_n5556_ = 1'b0;
endcase
casez ({new_n1421_, new_n5315_})
2'b01 : new_n5557_ = 1'b1;
default : new_n5557_ = 1'b0;
endcase
casez ({new_n559_, new_n5321_})
2'b01 : new_n5558_ = 1'b1;
default : new_n5558_ = 1'b0;
endcase
casez ({new_n3794_, new_n5337_})
2'b01 : new_n5559_ = 1'b1;
default : new_n5559_ = 1'b0;
endcase
casez ({new_n4748_, new_n5350_})
2'b11 : new_n5560_ = 1'b1;
default : new_n5560_ = 1'b0;
endcase
casez ({new_n4621_, new_n5352_})
2'b01 : new_n5561_ = 1'b1;
default : new_n5561_ = 1'b0;
endcase
casez ({new_n415_, new_n5354_})
2'b01 : new_n5562_ = 1'b1;
default : new_n5562_ = 1'b0;
endcase
casez ({new_n2302_, new_n5355_})
2'b11 : new_n5563_ = 1'b1;
default : new_n5563_ = 1'b0;
endcase
casez ({new_n690_, new_n5361_})
2'b01 : new_n5564_ = 1'b1;
default : new_n5564_ = 1'b0;
endcase
casez ({new_n1415_, new_n5369_})
2'b01 : new_n5565_ = 1'b1;
default : new_n5565_ = 1'b0;
endcase
casez ({new_n529_, new_n1176_})
2'b00 : new_n5566_ = 1'b1;
default : new_n5566_ = 1'b0;
endcase
casez ({new_n466_, new_n5376_})
2'b01 : new_n5567_ = 1'b1;
default : new_n5567_ = 1'b0;
endcase
casez ({new_n1052_, new_n5385_})
2'b01 : new_n5568_ = 1'b1;
default : new_n5568_ = 1'b0;
endcase
casez ({new_n4021_, new_n5386_})
2'b01 : new_n5569_ = 1'b1;
default : new_n5569_ = 1'b0;
endcase
casez ({new_n684_, new_n5405_})
2'b01 : new_n5570_ = 1'b1;
default : new_n5570_ = 1'b0;
endcase
casez ({new_n3785_, new_n5411_})
2'b01 : new_n5571_ = 1'b1;
default : new_n5571_ = 1'b0;
endcase
casez ({new_n1696_, new_n5413_})
2'b01 : new_n5572_ = 1'b1;
default : new_n5572_ = 1'b0;
endcase
casez ({new_n415_, new_n5425_})
2'b01 : new_n5573_ = 1'b1;
default : new_n5573_ = 1'b0;
endcase
casez ({new_n1193_, new_n1992_})
2'b00 : new_n5574_ = 1'b1;
default : new_n5574_ = 1'b0;
endcase
casez ({new_n2006_, new_n2008_})
2'b00 : new_n5575_ = 1'b1;
default : new_n5575_ = 1'b0;
endcase
casez ({new_n1198_, new_n2027_})
2'b00 : new_n5576_ = 1'b1;
default : new_n5576_ = 1'b0;
endcase
casez ({new_n2026_, new_n2035_})
2'b00 : new_n5577_ = 1'b1;
default : new_n5577_ = 1'b0;
endcase
casez ({new_n740_, new_n802_})
2'b00 : new_n5578_ = 1'b1;
default : new_n5578_ = 1'b0;
endcase
casez ({new_n2036_, new_n2044_})
2'b00 : new_n5579_ = 1'b1;
default : new_n5579_ = 1'b0;
endcase
casez ({new_n5930_, new_n808_})
2'b1? : new_n5580_ = 1'b1;
2'b?1 : new_n5580_ = 1'b1;
default : new_n5580_ = 1'b0;
endcase
casez ({new_n1663_, new_n2059_})
2'b01 : new_n5581_ = 1'b1;
default : new_n5581_ = 1'b0;
endcase
casez ({new_n2038_, new_n2071_})
2'b00 : new_n5582_ = 1'b1;
default : new_n5582_ = 1'b0;
endcase
casez ({new_n1513_, new_n2075_})
2'b11 : new_n5583_ = 1'b1;
default : new_n5583_ = 1'b0;
endcase
casez ({new_n590_, new_n1206_})
2'b00 : new_n5584_ = 1'b1;
default : new_n5584_ = 1'b0;
endcase
casez ({new_n2029_, new_n2080_})
2'b00 : new_n5585_ = 1'b1;
default : new_n5585_ = 1'b0;
endcase
casez ({new_n2013_, new_n2082_})
2'b00 : new_n5586_ = 1'b1;
default : new_n5586_ = 1'b0;
endcase
casez ({new_n85_, new_n291_, new_n1214_})
3'b11? : new_n5587_ = 1'b1;
3'b??1 : new_n5587_ = 1'b1;
default : new_n5587_ = 1'b0;
endcase
casez ({new_n521_, new_n816_})
2'b00 : new_n5588_ = 1'b1;
default : new_n5588_ = 1'b0;
endcase
casez ({new_n198_, new_n936_, new_n917_})
3'b10? : new_n5589_ = 1'b1;
3'b??1 : new_n5589_ = 1'b1;
default : new_n5589_ = 1'b0;
endcase
casez ({new_n1524_, new_n2119_})
2'b00 : new_n5590_ = 1'b1;
default : new_n5590_ = 1'b0;
endcase
casez ({new_n475_, new_n839_})
2'b00 : new_n5591_ = 1'b1;
default : new_n5591_ = 1'b0;
endcase
casez ({new_n1681_, new_n2160_})
2'b00 : new_n5592_ = 1'b1;
default : new_n5592_ = 1'b0;
endcase
casez ({u[2], new_n458_, new_n2163_})
3'b11? : new_n5593_ = 1'b1;
3'b??0 : new_n5593_ = 1'b1;
default : new_n5593_ = 1'b0;
endcase
casez ({new_n962_, new_n2166_})
2'b01 : new_n5594_ = 1'b1;
default : new_n5594_ = 1'b0;
endcase
casez ({new_n1326_, new_n2179_})
2'b01 : new_n5595_ = 1'b1;
default : new_n5595_ = 1'b0;
endcase
casez ({new_n617_, new_n1243_})
2'b00 : new_n5596_ = 1'b1;
default : new_n5596_ = 1'b0;
endcase
casez ({new_n687_, new_n853_})
2'b00 : new_n5597_ = 1'b1;
default : new_n5597_ = 1'b0;
endcase
casez ({new_n985_, new_n1243_})
2'b00 : new_n5598_ = 1'b1;
default : new_n5598_ = 1'b0;
endcase
casez ({new_n1017_, new_n2200_})
2'b01 : new_n5599_ = 1'b1;
default : new_n5599_ = 1'b0;
endcase
casez ({new_n410_, new_n553_})
2'b10 : new_n5600_ = 1'b1;
default : new_n5600_ = 1'b0;
endcase
casez ({new_n1841_, new_n2219_})
2'b01 : new_n5601_ = 1'b1;
default : new_n5601_ = 1'b0;
endcase
casez ({new_n207_, new_n263_, new_n560_})
3'b11? : new_n5602_ = 1'b1;
3'b??1 : new_n5602_ = 1'b1;
default : new_n5602_ = 1'b0;
endcase
casez ({new_n807_, new_n2237_})
2'b01 : new_n5603_ = 1'b1;
default : new_n5603_ = 1'b0;
endcase
casez ({new_n1745_, new_n2243_})
2'b01 : new_n5604_ = 1'b1;
default : new_n5604_ = 1'b0;
endcase
casez ({new_n917_, new_n1275_})
2'b00 : new_n5605_ = 1'b1;
default : new_n5605_ = 1'b0;
endcase
casez ({new_n560_, new_n563_})
2'b00 : new_n5606_ = 1'b1;
default : new_n5606_ = 1'b0;
endcase
casez ({new_n747_, new_n2260_})
2'b01 : new_n5607_ = 1'b1;
default : new_n5607_ = 1'b0;
endcase
casez ({new_n685_, new_n2265_})
2'b01 : new_n5608_ = 1'b1;
default : new_n5608_ = 1'b0;
endcase
casez ({new_n1693_, new_n2265_})
2'b01 : new_n5609_ = 1'b1;
default : new_n5609_ = 1'b0;
endcase
casez ({new_n1879_, new_n2273_})
2'b01 : new_n5610_ = 1'b1;
default : new_n5610_ = 1'b0;
endcase
casez ({new_n210_, new_n923_, new_n2277_})
3'b11? : new_n5611_ = 1'b1;
3'b??0 : new_n5611_ = 1'b1;
default : new_n5611_ = 1'b0;
endcase
casez ({new_n283_, new_n2287_})
2'b01 : new_n5612_ = 1'b1;
default : new_n5612_ = 1'b0;
endcase
casez ({new_n1893_, new_n2292_})
2'b01 : new_n5613_ = 1'b1;
default : new_n5613_ = 1'b0;
endcase
casez ({new_n550_, new_n2292_})
2'b11 : new_n5614_ = 1'b1;
default : new_n5614_ = 1'b0;
endcase
casez ({new_n759_, new_n1324_})
2'b10 : new_n5615_ = 1'b1;
default : new_n5615_ = 1'b0;
endcase
casez ({new_n1050_, new_n2304_})
2'b01 : new_n5616_ = 1'b1;
default : new_n5616_ = 1'b0;
endcase
casez ({new_n1590_, new_n2312_})
2'b01 : new_n5617_ = 1'b1;
default : new_n5617_ = 1'b0;
endcase
casez ({new_n562_, new_n2318_})
2'b01 : new_n5618_ = 1'b1;
default : new_n5618_ = 1'b0;
endcase
casez ({new_n1573_, new_n2326_})
2'b01 : new_n5619_ = 1'b1;
default : new_n5619_ = 1'b0;
endcase
casez ({new_n1697_, new_n2328_})
2'b01 : new_n5620_ = 1'b1;
default : new_n5620_ = 1'b0;
endcase
casez ({new_n83_, new_n396_, new_n2328_})
3'b11? : new_n5621_ = 1'b1;
3'b??0 : new_n5621_ = 1'b1;
default : new_n5621_ = 1'b0;
endcase
casez ({new_n521_, new_n1341_})
2'b00 : new_n5622_ = 1'b1;
default : new_n5622_ = 1'b0;
endcase
casez ({new_n642_, new_n2335_})
2'b00 : new_n5623_ = 1'b1;
default : new_n5623_ = 1'b0;
endcase
casez ({new_n1416_, new_n2335_})
2'b00 : new_n5624_ = 1'b1;
default : new_n5624_ = 1'b0;
endcase
casez ({new_n1555_, new_n2336_})
2'b00 : new_n5625_ = 1'b1;
default : new_n5625_ = 1'b0;
endcase
casez ({new_n562_, new_n1347_})
2'b00 : new_n5626_ = 1'b1;
default : new_n5626_ = 1'b0;
endcase
casez ({new_n419_, new_n890_})
2'b00 : new_n5627_ = 1'b1;
default : new_n5627_ = 1'b0;
endcase
casez ({new_n745_, new_n894_})
2'b00 : new_n5628_ = 1'b1;
default : new_n5628_ = 1'b0;
endcase
casez ({new_n562_, new_n896_})
2'b00 : new_n5629_ = 1'b1;
default : new_n5629_ = 1'b0;
endcase
casez ({new_n96_, new_n310_, new_n590_})
3'b01? : new_n5630_ = 1'b1;
3'b??1 : new_n5630_ = 1'b1;
default : new_n5630_ = 1'b0;
endcase
casez ({new_n232_, new_n311_})
2'b00 : new_n5631_ = 1'b1;
default : new_n5631_ = 1'b0;
endcase
casez ({new_n1243_, new_n1374_})
2'b00 : new_n5632_ = 1'b1;
default : new_n5632_ = 1'b0;
endcase
casez ({new_n670_, new_n1383_})
2'b00 : new_n5633_ = 1'b1;
default : new_n5633_ = 1'b0;
endcase
casez ({new_n760_, new_n909_})
2'b00 : new_n5634_ = 1'b1;
default : new_n5634_ = 1'b0;
endcase
casez ({new_n989_, new_n2507_})
2'b10 : new_n5635_ = 1'b1;
default : new_n5635_ = 1'b0;
endcase
casez ({new_n691_, new_n915_})
2'b00 : new_n5636_ = 1'b1;
default : new_n5636_ = 1'b0;
endcase
casez ({new_n833_, new_n915_})
2'b00 : new_n5637_ = 1'b1;
default : new_n5637_ = 1'b0;
endcase
casez ({new_n881_, new_n2564_})
2'b00 : new_n5638_ = 1'b1;
default : new_n5638_ = 1'b0;
endcase
casez ({new_n1360_, new_n1406_})
2'b00 : new_n5639_ = 1'b1;
default : new_n5639_ = 1'b0;
endcase
casez ({new_n782_, new_n1408_})
2'b00 : new_n5640_ = 1'b1;
default : new_n5640_ = 1'b0;
endcase
casez ({new_n1306_, new_n1410_})
2'b00 : new_n5641_ = 1'b1;
default : new_n5641_ = 1'b0;
endcase
casez ({new_n1313_, new_n1414_})
2'b00 : new_n5642_ = 1'b1;
default : new_n5642_ = 1'b0;
endcase
casez ({new_n577_, new_n1416_})
2'b00 : new_n5643_ = 1'b1;
default : new_n5643_ = 1'b0;
endcase
casez ({new_n973_, new_n1417_})
2'b00 : new_n5644_ = 1'b1;
default : new_n5644_ = 1'b0;
endcase
casez ({new_n645_, new_n1422_})
2'b00 : new_n5645_ = 1'b1;
default : new_n5645_ = 1'b0;
endcase
casez ({new_n232_, new_n618_})
2'b00 : new_n5646_ = 1'b1;
default : new_n5646_ = 1'b0;
endcase
casez ({new_n593_, new_n1427_})
2'b00 : new_n5647_ = 1'b1;
default : new_n5647_ = 1'b0;
endcase
casez ({new_n259_, new_n621_})
2'b00 : new_n5648_ = 1'b1;
default : new_n5648_ = 1'b0;
endcase
casez ({new_n2301_, new_n2630_})
2'b10 : new_n5649_ = 1'b1;
default : new_n5649_ = 1'b0;
endcase
casez ({new_n2261_, new_n2644_})
2'b10 : new_n5650_ = 1'b1;
default : new_n5650_ = 1'b0;
endcase
casez ({new_n1436_, new_n2644_})
2'b00 : new_n5651_ = 1'b1;
default : new_n5651_ = 1'b0;
endcase
casez ({new_n1048_, new_n2647_})
2'b00 : new_n5652_ = 1'b1;
default : new_n5652_ = 1'b0;
endcase
casez ({new_n1520_, new_n2648_})
2'b10 : new_n5653_ = 1'b1;
default : new_n5653_ = 1'b0;
endcase
casez ({new_n691_, new_n942_})
2'b00 : new_n5654_ = 1'b1;
default : new_n5654_ = 1'b0;
endcase
casez ({new_n521_, new_n2651_})
2'b00 : new_n5655_ = 1'b1;
default : new_n5655_ = 1'b0;
endcase
casez ({new_n1437_, new_n2668_})
2'b00 : new_n5656_ = 1'b1;
default : new_n5656_ = 1'b0;
endcase
casez ({new_n692_, new_n2671_})
2'b00 : new_n5657_ = 1'b1;
default : new_n5657_ = 1'b0;
endcase
casez ({new_n1407_, new_n2692_})
2'b00 : new_n5658_ = 1'b1;
default : new_n5658_ = 1'b0;
endcase
casez ({new_n1242_, new_n1469_})
2'b00 : new_n5659_ = 1'b1;
default : new_n5659_ = 1'b0;
endcase
casez ({new_n518_, new_n1469_})
2'b00 : new_n5660_ = 1'b1;
default : new_n5660_ = 1'b0;
endcase
casez ({new_n475_, new_n2713_})
2'b00 : new_n5661_ = 1'b1;
default : new_n5661_ = 1'b0;
endcase
casez ({new_n1696_, new_n2718_})
2'b00 : new_n5662_ = 1'b1;
default : new_n5662_ = 1'b0;
endcase
casez ({new_n704_, new_n2724_})
2'b00 : new_n5663_ = 1'b1;
default : new_n5663_ = 1'b0;
endcase
casez ({new_n1524_, new_n2727_})
2'b00 : new_n5664_ = 1'b1;
default : new_n5664_ = 1'b0;
endcase
casez ({new_n2336_, new_n2750_})
2'b00 : new_n5665_ = 1'b1;
default : new_n5665_ = 1'b0;
endcase
casez ({new_n1661_, new_n2760_})
2'b00 : new_n5666_ = 1'b1;
default : new_n5666_ = 1'b0;
endcase
casez ({new_n521_, new_n643_})
2'b00 : new_n5667_ = 1'b1;
default : new_n5667_ = 1'b0;
endcase
casez ({new_n504_, new_n967_})
2'b00 : new_n5668_ = 1'b1;
default : new_n5668_ = 1'b0;
endcase
casez ({new_n689_, new_n1497_})
2'b00 : new_n5669_ = 1'b1;
default : new_n5669_ = 1'b0;
endcase
casez ({new_n670_, new_n1498_})
2'b00 : new_n5670_ = 1'b1;
default : new_n5670_ = 1'b0;
endcase
casez ({new_n468_, new_n2806_})
2'b00 : new_n5671_ = 1'b1;
default : new_n5671_ = 1'b0;
endcase
casez ({new_n402_, new_n1513_})
2'b01 : new_n5672_ = 1'b1;
default : new_n5672_ = 1'b0;
endcase
casez ({new_n892_, new_n2833_})
2'b00 : new_n5673_ = 1'b1;
default : new_n5673_ = 1'b0;
endcase
casez ({new_n1055_, new_n1516_})
2'b01 : new_n5674_ = 1'b1;
default : new_n5674_ = 1'b0;
endcase
casez ({new_n1975_, new_n2844_})
2'b00 : new_n5675_ = 1'b1;
default : new_n5675_ = 1'b0;
endcase
casez ({new_n1436_, new_n1523_})
2'b00 : new_n5676_ = 1'b1;
default : new_n5676_ = 1'b0;
endcase
casez ({new_n807_, new_n1525_})
2'b00 : new_n5677_ = 1'b1;
default : new_n5677_ = 1'b0;
endcase
casez ({new_n286_, new_n650_})
2'b01 : new_n5678_ = 1'b1;
default : new_n5678_ = 1'b0;
endcase
casez ({new_n387_, new_n653_})
2'b00 : new_n5679_ = 1'b1;
default : new_n5679_ = 1'b0;
endcase
casez ({new_n1427_, new_n1571_})
2'b00 : new_n5680_ = 1'b1;
default : new_n5680_ = 1'b0;
endcase
casez ({new_n559_, new_n3100_})
2'b00 : new_n5681_ = 1'b1;
default : new_n5681_ = 1'b0;
endcase
casez ({new_n276_, new_n676_})
2'b00 : new_n5682_ = 1'b1;
default : new_n5682_ = 1'b0;
endcase
casez ({new_n802_, new_n1590_})
2'b00 : new_n5683_ = 1'b1;
default : new_n5683_ = 1'b0;
endcase
casez ({new_n1653_, new_n3157_})
2'b00 : new_n5684_ = 1'b1;
default : new_n5684_ = 1'b0;
endcase
casez ({new_n563_, new_n3160_})
2'b00 : new_n5685_ = 1'b1;
default : new_n5685_ = 1'b0;
endcase
casez ({new_n916_, new_n1594_})
2'b00 : new_n5686_ = 1'b1;
default : new_n5686_ = 1'b0;
endcase
casez ({new_n559_, new_n1597_})
2'b00 : new_n5687_ = 1'b1;
default : new_n5687_ = 1'b0;
endcase
casez ({new_n276_, new_n3196_})
2'b00 : new_n5688_ = 1'b1;
default : new_n5688_ = 1'b0;
endcase
casez ({new_n1693_, new_n3209_})
2'b00 : new_n5689_ = 1'b1;
default : new_n5689_ = 1'b0;
endcase
casez ({new_n759_, new_n1609_})
2'b10 : new_n5690_ = 1'b1;
default : new_n5690_ = 1'b0;
endcase
casez ({new_n565_, new_n686_})
2'b00 : new_n5691_ = 1'b1;
default : new_n5691_ = 1'b0;
endcase
casez ({new_n104_, new_n1025_, new_n546_})
3'b11? : new_n5692_ = 1'b1;
3'b??1 : new_n5692_ = 1'b1;
default : new_n5692_ = 1'b0;
endcase
casez ({new_n592_, new_n3338_})
2'b00 : new_n5693_ = 1'b1;
default : new_n5693_ = 1'b0;
endcase
casez ({new_n1664_, new_n3344_})
2'b00 : new_n5694_ = 1'b1;
default : new_n5694_ = 1'b0;
endcase
casez ({new_n609_, new_n3346_})
2'b00 : new_n5695_ = 1'b1;
default : new_n5695_ = 1'b0;
endcase
casez ({new_n2259_, new_n3349_})
2'b10 : new_n5696_ = 1'b1;
default : new_n5696_ = 1'b0;
endcase
casez ({new_n650_, new_n1626_})
2'b10 : new_n5697_ = 1'b1;
default : new_n5697_ = 1'b0;
endcase
casez ({new_n562_, new_n3413_})
2'b00 : new_n5698_ = 1'b1;
default : new_n5698_ = 1'b0;
endcase
casez ({new_n878_, new_n3439_})
2'b00 : new_n5699_ = 1'b1;
default : new_n5699_ = 1'b0;
endcase
casez ({new_n2301_, new_n3467_})
2'b10 : new_n5700_ = 1'b1;
default : new_n5700_ = 1'b0;
endcase
casez ({new_n609_, new_n3495_})
2'b00 : new_n5701_ = 1'b1;
default : new_n5701_ = 1'b0;
endcase
casez ({new_n461_, new_n1042_})
2'b00 : new_n5702_ = 1'b1;
default : new_n5702_ = 1'b0;
endcase
casez ({new_n368_, new_n703_})
2'b00 : new_n5703_ = 1'b1;
default : new_n5703_ = 1'b0;
endcase
casez ({new_n1109_, new_n1653_})
2'b00 : new_n5704_ = 1'b1;
default : new_n5704_ = 1'b0;
endcase
casez ({new_n326_, new_n3559_})
2'b00 : new_n5705_ = 1'b1;
default : new_n5705_ = 1'b0;
endcase
casez ({new_n811_, new_n1654_})
2'b00 : new_n5706_ = 1'b1;
default : new_n5706_ = 1'b0;
endcase
casez ({new_n409_, new_n704_})
2'b10 : new_n5707_ = 1'b1;
default : new_n5707_ = 1'b0;
endcase
casez ({new_n1310_, new_n1659_})
2'b00 : new_n5708_ = 1'b1;
default : new_n5708_ = 1'b0;
endcase
casez ({new_n584_, new_n1660_})
2'b00 : new_n5709_ = 1'b1;
default : new_n5709_ = 1'b0;
endcase
casez ({new_n506_, new_n1664_})
2'b00 : new_n5710_ = 1'b1;
default : new_n5710_ = 1'b0;
endcase
casez ({new_n723_, new_n1673_})
2'b00 : new_n5711_ = 1'b1;
default : new_n5711_ = 1'b0;
endcase
casez ({new_n975_, new_n1673_})
2'b00 : new_n5712_ = 1'b1;
default : new_n5712_ = 1'b0;
endcase
casez ({new_n1354_, new_n1674_})
2'b00 : new_n5713_ = 1'b1;
default : new_n5713_ = 1'b0;
endcase
casez ({new_n1417_, new_n3611_})
2'b00 : new_n5714_ = 1'b1;
default : new_n5714_ = 1'b0;
endcase
casez ({new_n690_, new_n1676_})
2'b00 : new_n5715_ = 1'b1;
default : new_n5715_ = 1'b0;
endcase
casez ({new_n1392_, new_n1678_})
2'b00 : new_n5716_ = 1'b1;
default : new_n5716_ = 1'b0;
endcase
casez ({new_n3302_, new_n3618_})
2'b00 : new_n5717_ = 1'b1;
default : new_n5717_ = 1'b0;
endcase
casez ({new_n297_, new_n1679_})
2'b00 : new_n5718_ = 1'b1;
default : new_n5718_ = 1'b0;
endcase
casez ({new_n983_, new_n3623_})
2'b00 : new_n5719_ = 1'b1;
default : new_n5719_ = 1'b0;
endcase
casez ({new_n653_, new_n3625_})
2'b00 : new_n5720_ = 1'b1;
default : new_n5720_ = 1'b0;
endcase
casez ({new_n827_, new_n1682_})
2'b00 : new_n5721_ = 1'b1;
default : new_n5721_ = 1'b0;
endcase
casez ({new_n1495_, new_n1684_})
2'b00 : new_n5722_ = 1'b1;
default : new_n5722_ = 1'b0;
endcase
casez ({new_n128_, new_n1686_})
2'b00 : new_n5723_ = 1'b1;
default : new_n5723_ = 1'b0;
endcase
casez ({new_n1584_, new_n3650_})
2'b00 : new_n5724_ = 1'b1;
default : new_n5724_ = 1'b0;
endcase
casez ({new_n2840_, new_n3651_})
2'b00 : new_n5725_ = 1'b1;
default : new_n5725_ = 1'b0;
endcase
casez ({new_n866_, new_n1689_})
2'b00 : new_n5726_ = 1'b1;
default : new_n5726_ = 1'b0;
endcase
casez ({new_n717_, new_n3654_})
2'b00 : new_n5727_ = 1'b1;
default : new_n5727_ = 1'b0;
endcase
casez ({new_n1499_, new_n1690_})
2'b00 : new_n5728_ = 1'b1;
default : new_n5728_ = 1'b0;
endcase
casez ({new_n2837_, new_n3657_})
2'b00 : new_n5729_ = 1'b1;
default : new_n5729_ = 1'b0;
endcase
casez ({new_n1730_, new_n3659_})
2'b00 : new_n5730_ = 1'b1;
default : new_n5730_ = 1'b0;
endcase
casez ({new_n2685_, new_n3664_})
2'b00 : new_n5731_ = 1'b1;
default : new_n5731_ = 1'b0;
endcase
casez ({new_n1862_, new_n3665_})
2'b00 : new_n5732_ = 1'b1;
default : new_n5732_ = 1'b0;
endcase
casez ({new_n1480_, new_n1694_})
2'b00 : new_n5733_ = 1'b1;
default : new_n5733_ = 1'b0;
endcase
casez ({new_n521_, new_n1056_})
2'b00 : new_n5734_ = 1'b1;
default : new_n5734_ = 1'b0;
endcase
casez ({new_n1199_, new_n3674_})
2'b00 : new_n5735_ = 1'b1;
default : new_n5735_ = 1'b0;
endcase
casez ({new_n1840_, new_n3677_})
2'b00 : new_n5736_ = 1'b1;
default : new_n5736_ = 1'b0;
endcase
casez ({new_n1665_, new_n1697_})
2'b00 : new_n5737_ = 1'b1;
default : new_n5737_ = 1'b0;
endcase
casez ({new_n1585_, new_n3692_})
2'b00 : new_n5738_ = 1'b1;
default : new_n5738_ = 1'b0;
endcase
casez ({new_n468_, new_n1060_})
2'b00 : new_n5739_ = 1'b1;
default : new_n5739_ = 1'b0;
endcase
casez ({new_n1660_, new_n3739_})
2'b01 : new_n5740_ = 1'b1;
default : new_n5740_ = 1'b0;
endcase
casez ({new_n474_, new_n1715_})
2'b00 : new_n5741_ = 1'b1;
default : new_n5741_ = 1'b0;
endcase
casez ({new_n2697_, new_n3742_})
2'b00 : new_n5742_ = 1'b1;
default : new_n5742_ = 1'b0;
endcase
casez ({new_n1603_, new_n3743_})
2'b00 : new_n5743_ = 1'b1;
default : new_n5743_ = 1'b0;
endcase
casez ({new_n1031_, new_n3752_})
2'b00 : new_n5744_ = 1'b1;
default : new_n5744_ = 1'b0;
endcase
casez ({new_n3427_, new_n3757_})
2'b00 : new_n5745_ = 1'b1;
default : new_n5745_ = 1'b0;
endcase
casez ({new_n583_, new_n3763_})
2'b00 : new_n5746_ = 1'b1;
default : new_n5746_ = 1'b0;
endcase
casez ({new_n765_, new_n800_, new_n3784_})
3'b11? : new_n5747_ = 1'b1;
3'b??1 : new_n5747_ = 1'b1;
default : new_n5747_ = 1'b0;
endcase
casez ({new_n907_, new_n3788_})
2'b00 : new_n5748_ = 1'b1;
default : new_n5748_ = 1'b0;
endcase
casez ({new_n1227_, new_n3793_})
2'b00 : new_n5749_ = 1'b1;
default : new_n5749_ = 1'b0;
endcase
casez ({new_n813_, new_n3812_})
2'b00 : new_n5750_ = 1'b1;
default : new_n5750_ = 1'b0;
endcase
casez ({new_n233_, new_n3813_})
2'b00 : new_n5751_ = 1'b1;
default : new_n5751_ = 1'b0;
endcase
casez ({new_n1464_, new_n3819_})
2'b00 : new_n5752_ = 1'b1;
default : new_n5752_ = 1'b0;
endcase
casez ({new_n1666_, new_n1727_})
2'b00 : new_n5753_ = 1'b1;
default : new_n5753_ = 1'b0;
endcase
casez ({new_n1593_, new_n3830_})
2'b00 : new_n5754_ = 1'b1;
default : new_n5754_ = 1'b0;
endcase
casez ({new_n2799_, new_n3834_})
2'b00 : new_n5755_ = 1'b1;
default : new_n5755_ = 1'b0;
endcase
casez ({new_n547_, new_n3837_})
2'b00 : new_n5756_ = 1'b1;
default : new_n5756_ = 1'b0;
endcase
casez ({new_n3131_, new_n3844_})
2'b10 : new_n5757_ = 1'b1;
default : new_n5757_ = 1'b0;
endcase
casez ({new_n470_, new_n3857_})
2'b00 : new_n5758_ = 1'b1;
default : new_n5758_ = 1'b0;
endcase
casez ({new_n2795_, new_n3861_})
2'b00 : new_n5759_ = 1'b1;
default : new_n5759_ = 1'b0;
endcase
casez ({new_n896_, new_n3877_})
2'b01 : new_n5760_ = 1'b1;
default : new_n5760_ = 1'b0;
endcase
casez ({new_n1897_, new_n3879_})
2'b00 : new_n5761_ = 1'b1;
default : new_n5761_ = 1'b0;
endcase
casez ({new_n811_, new_n3882_})
2'b00 : new_n5762_ = 1'b1;
default : new_n5762_ = 1'b0;
endcase
casez ({new_n758_, new_n1734_})
2'b10 : new_n5763_ = 1'b1;
default : new_n5763_ = 1'b0;
endcase
casez ({new_n2797_, new_n3887_})
2'b00 : new_n5764_ = 1'b1;
default : new_n5764_ = 1'b0;
endcase
casez ({new_n1133_, new_n3890_})
2'b00 : new_n5765_ = 1'b1;
default : new_n5765_ = 1'b0;
endcase
casez ({new_n3341_, new_n3903_})
2'b00 : new_n5766_ = 1'b1;
default : new_n5766_ = 1'b0;
endcase
casez ({new_n3798_, new_n3906_})
2'b01 : new_n5767_ = 1'b1;
default : new_n5767_ = 1'b0;
endcase
casez ({new_n895_, new_n1070_})
2'b00 : new_n5768_ = 1'b1;
default : new_n5768_ = 1'b0;
endcase
casez ({new_n1066_, new_n3910_})
2'b00 : new_n5769_ = 1'b1;
default : new_n5769_ = 1'b0;
endcase
casez ({new_n1642_, new_n3917_})
2'b00 : new_n5770_ = 1'b1;
default : new_n5770_ = 1'b0;
endcase
casez ({new_n1066_, new_n3918_})
2'b00 : new_n5771_ = 1'b1;
default : new_n5771_ = 1'b0;
endcase
casez ({new_n806_, new_n1739_})
2'b00 : new_n5772_ = 1'b1;
default : new_n5772_ = 1'b0;
endcase
casez ({new_n1615_, new_n3923_})
2'b00 : new_n5773_ = 1'b1;
default : new_n5773_ = 1'b0;
endcase
casez ({new_n1604_, new_n3930_})
2'b00 : new_n5774_ = 1'b1;
default : new_n5774_ = 1'b0;
endcase
casez ({new_n587_, new_n3939_})
2'b00 : new_n5775_ = 1'b1;
default : new_n5775_ = 1'b0;
endcase
casez ({new_n178_, new_n712_, new_n3940_})
3'b11? : new_n5776_ = 1'b1;
3'b??1 : new_n5776_ = 1'b1;
default : new_n5776_ = 1'b0;
endcase
casez ({new_n1124_, new_n3942_})
2'b00 : new_n5777_ = 1'b1;
default : new_n5777_ = 1'b0;
endcase
casez ({u[1], new_n2781_, new_n3947_})
3'b11? : new_n5778_ = 1'b1;
3'b??1 : new_n5778_ = 1'b1;
default : new_n5778_ = 1'b0;
endcase
casez ({new_n3669_, new_n3951_})
2'b00 : new_n5779_ = 1'b1;
default : new_n5779_ = 1'b0;
endcase
casez ({new_n373_, new_n3950_})
2'b00 : new_n5780_ = 1'b1;
default : new_n5780_ = 1'b0;
endcase
casez ({new_n292_, new_n3963_})
2'b00 : new_n5781_ = 1'b1;
default : new_n5781_ = 1'b0;
endcase
casez ({new_n1837_, new_n3965_})
2'b00 : new_n5782_ = 1'b1;
default : new_n5782_ = 1'b0;
endcase
casez ({new_n461_, new_n3969_})
2'b01 : new_n5783_ = 1'b1;
default : new_n5783_ = 1'b0;
endcase
casez ({new_n1072_, new_n3970_})
2'b00 : new_n5784_ = 1'b1;
default : new_n5784_ = 1'b0;
endcase
casez ({new_n3850_, new_n3974_})
2'b01 : new_n5785_ = 1'b1;
default : new_n5785_ = 1'b0;
endcase
casez ({new_n2334_, new_n3982_})
2'b01 : new_n5786_ = 1'b1;
default : new_n5786_ = 1'b0;
endcase
casez ({new_n2995_, new_n3999_})
2'b00 : new_n5787_ = 1'b1;
default : new_n5787_ = 1'b0;
endcase
casez ({new_n3797_, new_n4001_})
2'b01 : new_n5788_ = 1'b1;
default : new_n5788_ = 1'b0;
endcase
casez ({new_n1415_, new_n4010_})
2'b00 : new_n5789_ = 1'b1;
default : new_n5789_ = 1'b0;
endcase
casez ({new_n326_, new_n1753_})
2'b00 : new_n5790_ = 1'b1;
default : new_n5790_ = 1'b0;
endcase
casez ({new_n1487_, new_n4044_})
2'b00 : new_n5791_ = 1'b1;
default : new_n5791_ = 1'b0;
endcase
casez ({new_n245_, new_n1087_})
2'b00 : new_n5792_ = 1'b1;
default : new_n5792_ = 1'b0;
endcase
casez ({new_n885_, new_n4053_})
2'b00 : new_n5793_ = 1'b1;
default : new_n5793_ = 1'b0;
endcase
casez ({new_n450_, new_n1087_})
2'b00 : new_n5794_ = 1'b1;
default : new_n5794_ = 1'b0;
endcase
casez ({new_n972_, new_n1087_})
2'b10 : new_n5795_ = 1'b1;
default : new_n5795_ = 1'b0;
endcase
casez ({new_n2287_, new_n4060_})
2'b11 : new_n5796_ = 1'b1;
default : new_n5796_ = 1'b0;
endcase
casez ({new_n590_, new_n4063_})
2'b00 : new_n5797_ = 1'b1;
default : new_n5797_ = 1'b0;
endcase
casez ({new_n92_, new_n1765_, new_n847_})
3'b10? : new_n5798_ = 1'b1;
3'b??1 : new_n5798_ = 1'b1;
default : new_n5798_ = 1'b0;
endcase
casez ({new_n2273_, new_n4064_})
2'b11 : new_n5799_ = 1'b1;
default : new_n5799_ = 1'b0;
endcase
casez ({new_n1735_, new_n4071_})
2'b00 : new_n5800_ = 1'b1;
default : new_n5800_ = 1'b0;
endcase
casez ({new_n2028_, new_n4076_})
2'b10 : new_n5801_ = 1'b1;
default : new_n5801_ = 1'b0;
endcase
casez ({new_n2111_, new_n4087_})
2'b00 : new_n5802_ = 1'b1;
default : new_n5802_ = 1'b0;
endcase
casez ({new_n2807_, new_n4092_})
2'b00 : new_n5803_ = 1'b1;
default : new_n5803_ = 1'b0;
endcase
casez ({new_n3978_, new_n4091_})
2'b01 : new_n5804_ = 1'b1;
default : new_n5804_ = 1'b0;
endcase
casez ({new_n3289_, new_n4103_})
2'b00 : new_n5805_ = 1'b1;
default : new_n5805_ = 1'b0;
endcase
casez ({new_n1681_, new_n4110_})
2'b01 : new_n5806_ = 1'b1;
default : new_n5806_ = 1'b0;
endcase
casez ({new_n1472_, new_n4114_})
2'b00 : new_n5807_ = 1'b1;
default : new_n5807_ = 1'b0;
endcase
casez ({new_n488_, new_n1096_, new_n547_})
3'b11? : new_n5808_ = 1'b1;
3'b??1 : new_n5808_ = 1'b1;
default : new_n5808_ = 1'b0;
endcase
casez ({new_n1471_, new_n4121_})
2'b00 : new_n5809_ = 1'b1;
default : new_n5809_ = 1'b0;
endcase
casez ({new_n698_, new_n4129_})
2'b00 : new_n5810_ = 1'b1;
default : new_n5810_ = 1'b0;
endcase
casez ({new_n1705_, new_n4164_})
2'b01 : new_n5811_ = 1'b1;
default : new_n5811_ = 1'b0;
endcase
casez ({new_n653_, new_n1099_})
2'b00 : new_n5812_ = 1'b1;
default : new_n5812_ = 1'b0;
endcase
casez ({new_n1875_, new_n4173_})
2'b00 : new_n5813_ = 1'b1;
default : new_n5813_ = 1'b0;
endcase
casez ({new_n1191_, new_n4174_})
2'b10 : new_n5814_ = 1'b1;
default : new_n5814_ = 1'b0;
endcase
casez ({new_n1692_, new_n4177_})
2'b00 : new_n5815_ = 1'b1;
default : new_n5815_ = 1'b0;
endcase
casez ({new_n826_, new_n4188_})
2'b00 : new_n5816_ = 1'b1;
default : new_n5816_ = 1'b0;
endcase
casez ({new_n3886_, new_n4183_})
2'b01 : new_n5817_ = 1'b1;
default : new_n5817_ = 1'b0;
endcase
casez ({new_n415_, new_n4191_})
2'b01 : new_n5818_ = 1'b1;
default : new_n5818_ = 1'b0;
endcase
casez ({new_n1884_, new_n4192_})
2'b00 : new_n5819_ = 1'b1;
default : new_n5819_ = 1'b0;
endcase
casez ({new_n429_, new_n4220_})
2'b00 : new_n5820_ = 1'b1;
default : new_n5820_ = 1'b0;
endcase
casez ({new_n1675_, new_n4233_})
2'b00 : new_n5821_ = 1'b1;
default : new_n5821_ = 1'b0;
endcase
casez ({new_n2200_, new_n4236_})
2'b10 : new_n5822_ = 1'b1;
default : new_n5822_ = 1'b0;
endcase
casez ({new_n1299_, new_n4240_})
2'b00 : new_n5823_ = 1'b1;
default : new_n5823_ = 1'b0;
endcase
casez ({new_n1747_, new_n4247_})
2'b00 : new_n5824_ = 1'b1;
default : new_n5824_ = 1'b0;
endcase
casez ({new_n1523_, new_n4254_})
2'b00 : new_n5825_ = 1'b1;
default : new_n5825_ = 1'b0;
endcase
casez ({new_n1280_, new_n4255_})
2'b00 : new_n5826_ = 1'b1;
default : new_n5826_ = 1'b0;
endcase
casez ({new_n4014_, new_n4259_})
2'b01 : new_n5827_ = 1'b1;
default : new_n5827_ = 1'b0;
endcase
casez ({new_n1838_, new_n4262_})
2'b00 : new_n5828_ = 1'b1;
default : new_n5828_ = 1'b0;
endcase
casez ({new_n1836_, new_n4264_})
2'b00 : new_n5829_ = 1'b1;
default : new_n5829_ = 1'b0;
endcase
casez ({new_n519_, new_n4266_})
2'b00 : new_n5830_ = 1'b1;
default : new_n5830_ = 1'b0;
endcase
casez ({new_n1413_, new_n4269_})
2'b10 : new_n5831_ = 1'b1;
default : new_n5831_ = 1'b0;
endcase
casez ({new_n1751_, new_n4270_})
2'b00 : new_n5832_ = 1'b1;
default : new_n5832_ = 1'b0;
endcase
casez ({new_n3397_, new_n4273_})
2'b00 : new_n5833_ = 1'b1;
default : new_n5833_ = 1'b0;
endcase
casez ({new_n1691_, new_n4287_})
2'b00 : new_n5834_ = 1'b1;
default : new_n5834_ = 1'b0;
endcase
casez ({new_n3856_, new_n4301_})
2'b01 : new_n5835_ = 1'b1;
default : new_n5835_ = 1'b0;
endcase
casez ({new_n4100_, new_n4304_})
2'b10 : new_n5836_ = 1'b1;
default : new_n5836_ = 1'b0;
endcase
casez ({new_n3697_, new_n4308_})
2'b00 : new_n5837_ = 1'b1;
default : new_n5837_ = 1'b0;
endcase
casez ({new_n1855_, new_n4312_})
2'b00 : new_n5838_ = 1'b1;
default : new_n5838_ = 1'b0;
endcase
casez ({new_n1734_, new_n4313_})
2'b00 : new_n5839_ = 1'b1;
default : new_n5839_ = 1'b0;
endcase
casez ({new_n3059_, new_n4311_})
2'b00 : new_n5840_ = 1'b1;
default : new_n5840_ = 1'b0;
endcase
casez ({new_n2267_, new_n4316_})
2'b11 : new_n5841_ = 1'b1;
default : new_n5841_ = 1'b0;
endcase
casez ({new_n3885_, new_n4318_})
2'b10 : new_n5842_ = 1'b1;
default : new_n5842_ = 1'b0;
endcase
casez ({new_n1275_, new_n4323_})
2'b00 : new_n5843_ = 1'b1;
default : new_n5843_ = 1'b0;
endcase
casez ({new_n3769_, new_n4324_})
2'b01 : new_n5844_ = 1'b1;
default : new_n5844_ = 1'b0;
endcase
casez ({new_n1667_, new_n4329_})
2'b01 : new_n5845_ = 1'b1;
default : new_n5845_ = 1'b0;
endcase
casez ({new_n435_, new_n4337_})
2'b00 : new_n5846_ = 1'b1;
default : new_n5846_ = 1'b0;
endcase
casez ({new_n3620_, new_n4350_})
2'b01 : new_n5847_ = 1'b1;
default : new_n5847_ = 1'b0;
endcase
casez ({new_n3042_, new_n4364_})
2'b00 : new_n5848_ = 1'b1;
default : new_n5848_ = 1'b0;
endcase
casez ({new_n2846_, new_n4367_})
2'b00 : new_n5849_ = 1'b1;
default : new_n5849_ = 1'b0;
endcase
casez ({new_n1520_, new_n1829_})
2'b10 : new_n5850_ = 1'b1;
default : new_n5850_ = 1'b0;
endcase
casez ({new_n546_, new_n1832_})
2'b00 : new_n5851_ = 1'b1;
default : new_n5851_ = 1'b0;
endcase
casez ({new_n3737_, new_n4393_})
2'b01 : new_n5852_ = 1'b1;
default : new_n5852_ = 1'b0;
endcase
casez ({new_n3921_, new_n4395_})
2'b01 : new_n5853_ = 1'b1;
default : new_n5853_ = 1'b0;
endcase
casez ({new_n684_, new_n1837_})
2'b00 : new_n5854_ = 1'b1;
default : new_n5854_ = 1'b0;
endcase
casez ({new_n1682_, new_n4433_})
2'b00 : new_n5855_ = 1'b1;
default : new_n5855_ = 1'b0;
endcase
casez ({new_n107_, new_n456_, new_n4439_})
3'b01? : new_n5856_ = 1'b1;
3'b??1 : new_n5856_ = 1'b1;
default : new_n5856_ = 1'b0;
endcase
casez ({new_n1675_, new_n4440_})
2'b00 : new_n5857_ = 1'b1;
default : new_n5857_ = 1'b0;
endcase
casez ({new_n1408_, new_n4457_})
2'b00 : new_n5858_ = 1'b1;
default : new_n5858_ = 1'b0;
endcase
casez ({new_n320_, new_n435_, new_n4474_})
3'b01? : new_n5859_ = 1'b1;
3'b??1 : new_n5859_ = 1'b1;
default : new_n5859_ = 1'b0;
endcase
casez ({new_n904_, new_n4480_})
2'b00 : new_n5860_ = 1'b1;
default : new_n5860_ = 1'b0;
endcase
casez ({new_n3684_, new_n4485_})
2'b01 : new_n5861_ = 1'b1;
default : new_n5861_ = 1'b0;
endcase
casez ({new_n1689_, new_n4495_})
2'b00 : new_n5862_ = 1'b1;
default : new_n5862_ = 1'b0;
endcase
casez ({new_n1452_, new_n4505_})
2'b00 : new_n5863_ = 1'b1;
default : new_n5863_ = 1'b0;
endcase
casez ({new_n1502_, new_n4511_})
2'b00 : new_n5864_ = 1'b1;
default : new_n5864_ = 1'b0;
endcase
casez ({new_n1887_, new_n4514_})
2'b00 : new_n5865_ = 1'b1;
default : new_n5865_ = 1'b0;
endcase
casez ({new_n546_, new_n4515_})
2'b00 : new_n5866_ = 1'b1;
default : new_n5866_ = 1'b0;
endcase
casez ({new_n1749_, new_n4520_})
2'b00 : new_n5867_ = 1'b1;
default : new_n5867_ = 1'b0;
endcase
casez ({new_n2803_, new_n4525_})
2'b00 : new_n5868_ = 1'b1;
default : new_n5868_ = 1'b0;
endcase
casez ({new_n546_, new_n4536_})
2'b01 : new_n5869_ = 1'b1;
default : new_n5869_ = 1'b0;
endcase
casez ({new_n93_, new_n354_, new_n4540_})
3'b11? : new_n5870_ = 1'b1;
3'b??0 : new_n5870_ = 1'b1;
default : new_n5870_ = 1'b0;
endcase
casez ({x[1], new_n104_, new_n269_, new_n4552_})
4'b101? : new_n5871_ = 1'b1;
4'b???1 : new_n5871_ = 1'b1;
default : new_n5871_ = 1'b0;
endcase
casez ({new_n1692_, new_n4558_})
2'b00 : new_n5872_ = 1'b1;
default : new_n5872_ = 1'b0;
endcase
casez ({y[2], new_n197_, new_n4560_})
3'b01? : new_n5873_ = 1'b1;
3'b??1 : new_n5873_ = 1'b1;
default : new_n5873_ = 1'b0;
endcase
casez ({new_n3265_, new_n4569_})
2'b00 : new_n5874_ = 1'b1;
default : new_n5874_ = 1'b0;
endcase
casez ({new_n646_, new_n4571_})
2'b00 : new_n5875_ = 1'b1;
default : new_n5875_ = 1'b0;
endcase
casez ({new_n1654_, new_n1860_})
2'b00 : new_n5876_ = 1'b1;
default : new_n5876_ = 1'b0;
endcase
casez ({new_n1701_, new_n4617_})
2'b00 : new_n5877_ = 1'b1;
default : new_n5877_ = 1'b0;
endcase
casez ({new_n3128_, new_n4679_})
2'b01 : new_n5878_ = 1'b1;
default : new_n5878_ = 1'b0;
endcase
casez ({new_n2125_, new_n4680_})
2'b01 : new_n5879_ = 1'b1;
default : new_n5879_ = 1'b0;
endcase
casez ({new_n1481_, new_n4684_})
2'b01 : new_n5880_ = 1'b1;
default : new_n5880_ = 1'b0;
endcase
casez ({new_n3111_, new_n4693_})
2'b01 : new_n5881_ = 1'b1;
default : new_n5881_ = 1'b0;
endcase
casez ({new_n819_, new_n1876_})
2'b00 : new_n5882_ = 1'b1;
default : new_n5882_ = 1'b0;
endcase
casez ({new_n474_, new_n4697_})
2'b01 : new_n5883_ = 1'b1;
default : new_n5883_ = 1'b0;
endcase
casez ({new_n3959_, new_n4698_})
2'b11 : new_n5884_ = 1'b1;
default : new_n5884_ = 1'b0;
endcase
casez ({new_n1277_, new_n4702_})
2'b01 : new_n5885_ = 1'b1;
default : new_n5885_ = 1'b0;
endcase
casez ({new_n655_, new_n4704_})
2'b01 : new_n5886_ = 1'b1;
default : new_n5886_ = 1'b0;
endcase
casez ({new_n2840_, new_n4705_})
2'b01 : new_n5887_ = 1'b1;
default : new_n5887_ = 1'b0;
endcase
casez ({new_n1732_, new_n4706_})
2'b01 : new_n5888_ = 1'b1;
default : new_n5888_ = 1'b0;
endcase
casez ({new_n1453_, new_n4707_})
2'b01 : new_n5889_ = 1'b1;
default : new_n5889_ = 1'b0;
endcase
casez ({new_n4630_, new_n4708_})
2'b01 : new_n5890_ = 1'b1;
default : new_n5890_ = 1'b0;
endcase
casez ({new_n4494_, new_n4710_})
2'b01 : new_n5891_ = 1'b1;
default : new_n5891_ = 1'b0;
endcase
casez ({new_n645_, new_n759_})
2'b01 : new_n5892_ = 1'b1;
default : new_n5892_ = 1'b0;
endcase
casez ({new_n4054_, new_n4721_})
2'b11 : new_n5893_ = 1'b1;
default : new_n5893_ = 1'b0;
endcase
casez ({new_n1279_, new_n4723_})
2'b01 : new_n5894_ = 1'b1;
default : new_n5894_ = 1'b0;
endcase
casez ({new_n1139_, new_n4725_})
2'b01 : new_n5895_ = 1'b1;
default : new_n5895_ = 1'b0;
endcase
casez ({new_n1480_, new_n4734_})
2'b01 : new_n5896_ = 1'b1;
default : new_n5896_ = 1'b0;
endcase
casez ({new_n3632_, new_n4735_})
2'b01 : new_n5897_ = 1'b1;
default : new_n5897_ = 1'b0;
endcase
casez ({new_n2628_, new_n4736_})
2'b01 : new_n5898_ = 1'b1;
default : new_n5898_ = 1'b0;
endcase
casez ({new_n3252_, new_n4740_})
2'b01 : new_n5899_ = 1'b1;
default : new_n5899_ = 1'b0;
endcase
casez ({new_n1669_, new_n4751_})
2'b01 : new_n5900_ = 1'b1;
default : new_n5900_ = 1'b0;
endcase
casez ({new_n196_, new_n263_, new_n4756_})
3'b11? : new_n5901_ = 1'b1;
3'b??0 : new_n5901_ = 1'b1;
default : new_n5901_ = 1'b0;
endcase
casez ({new_n1728_, new_n4764_})
2'b01 : new_n5902_ = 1'b1;
default : new_n5902_ = 1'b0;
endcase
casez ({new_n4538_, new_n4769_})
2'b11 : new_n5903_ = 1'b1;
default : new_n5903_ = 1'b0;
endcase
casez ({new_n3046_, new_n4771_})
2'b01 : new_n5904_ = 1'b1;
default : new_n5904_ = 1'b0;
endcase
casez ({new_n2194_, new_n4778_})
2'b11 : new_n5905_ = 1'b1;
default : new_n5905_ = 1'b0;
endcase
casez ({new_n1730_, new_n4792_})
2'b01 : new_n5906_ = 1'b1;
default : new_n5906_ = 1'b0;
endcase
casez ({new_n4043_, new_n4793_})
2'b11 : new_n5907_ = 1'b1;
default : new_n5907_ = 1'b0;
endcase
casez ({new_n1837_, new_n4796_})
2'b01 : new_n5908_ = 1'b1;
default : new_n5908_ = 1'b0;
endcase
casez ({new_n4267_, new_n4797_})
2'b11 : new_n5909_ = 1'b1;
default : new_n5909_ = 1'b0;
endcase
casez ({new_n2684_, new_n4803_})
2'b01 : new_n5910_ = 1'b1;
default : new_n5910_ = 1'b0;
endcase
casez ({new_n3242_, new_n4809_})
2'b01 : new_n5911_ = 1'b1;
default : new_n5911_ = 1'b0;
endcase
casez ({new_n3765_, new_n4816_})
2'b01 : new_n5912_ = 1'b1;
default : new_n5912_ = 1'b0;
endcase
casez ({new_n4144_, new_n4822_})
2'b01 : new_n5913_ = 1'b1;
default : new_n5913_ = 1'b0;
endcase
casez ({new_n2692_, new_n4823_})
2'b01 : new_n5914_ = 1'b1;
default : new_n5914_ = 1'b0;
endcase
casez ({new_n1056_, new_n4826_})
2'b01 : new_n5915_ = 1'b1;
default : new_n5915_ = 1'b0;
endcase
casez ({new_n1852_, new_n4827_})
2'b01 : new_n5916_ = 1'b1;
default : new_n5916_ = 1'b0;
endcase
casez ({new_n2241_, new_n4833_})
2'b11 : new_n5917_ = 1'b1;
default : new_n5917_ = 1'b0;
endcase
casez ({new_n3916_, new_n4835_})
2'b01 : new_n5918_ = 1'b1;
default : new_n5918_ = 1'b0;
endcase
casez ({new_n759_, new_n4846_})
2'b11 : new_n5919_ = 1'b1;
default : new_n5919_ = 1'b0;
endcase
casez ({new_n184_, new_n819_})
2'b11 : new_n5920_ = 1'b1;
default : new_n5920_ = 1'b0;
endcase
casez ({new_n307_, new_n562_})
2'b11 : new_n5921_ = 1'b1;
default : new_n5921_ = 1'b0;
endcase
casez ({new_n396_, new_n563_})
2'b11 : new_n5922_ = 1'b1;
default : new_n5922_ = 1'b0;
endcase
casez ({new_n98_, new_n884_})
2'b11 : new_n5923_ = 1'b1;
default : new_n5923_ = 1'b0;
endcase
casez ({new_n121_, new_n588_})
2'b11 : new_n5924_ = 1'b1;
default : new_n5924_ = 1'b0;
endcase
casez ({new_n174_, new_n915_})
2'b11 : new_n5925_ = 1'b1;
default : new_n5925_ = 1'b0;
endcase
casez ({new_n87_, new_n1526_})
2'b11 : new_n5926_ = 1'b1;
default : new_n5926_ = 1'b0;
endcase
casez ({new_n517_, new_n653_})
2'b11 : new_n5927_ = 1'b1;
default : new_n5927_ = 1'b0;
endcase
casez ({new_n323_, new_n703_})
2'b11 : new_n5928_ = 1'b1;
default : new_n5928_ = 1'b0;
endcase
casez ({new_n109_, new_n232_})
2'b01 : new_n5929_ = 1'b1;
default : new_n5929_ = 1'b0;
endcase
casez ({new_n117_, new_n250_})
2'b11 : new_n5930_ = 1'b1;
default : new_n5930_ = 1'b0;
endcase
casez ({new_n2429_, new_n4859_})
2'b01 : new_n5931_ = 1'b1;
default : new_n5931_ = 1'b0;
endcase
casez ({new_n1719_, new_n4858_})
2'b00 : new_n5932_ = 1'b1;
default : new_n5932_ = 1'b0;
endcase
casez ({new_n1084_, new_n1918_})
2'b00 : new_n5933_ = 1'b1;
default : new_n5933_ = 1'b0;
endcase
casez ({new_n595_, new_n4854_})
2'b01 : new_n5934_ = 1'b1;
default : new_n5934_ = 1'b0;
endcase
casez ({new_n1489_, new_n4876_})
2'b00 : new_n5935_ = 1'b1;
default : new_n5935_ = 1'b0;
endcase
casez ({new_n2708_, new_n4875_})
2'b00 : new_n5936_ = 1'b1;
default : new_n5936_ = 1'b0;
endcase
casez ({new_n2335_, new_n4907_})
2'b00 : new_n5937_ = 1'b1;
default : new_n5937_ = 1'b0;
endcase
casez ({new_n1478_, new_n4928_})
2'b00 : new_n5938_ = 1'b1;
default : new_n5938_ = 1'b0;
endcase
casez ({new_n2337_, new_n4948_})
2'b11 : new_n5939_ = 1'b1;
default : new_n5939_ = 1'b0;
endcase
casez ({new_n4993_, new_n5003_})
2'b01 : new_n5940_ = 1'b1;
default : new_n5940_ = 1'b0;
endcase
casez ({new_n4766_, new_n5012_})
2'b10 : new_n5941_ = 1'b1;
default : new_n5941_ = 1'b0;
endcase
casez ({new_n4807_, new_n5023_})
2'b01 : new_n5942_ = 1'b1;
default : new_n5942_ = 1'b0;
endcase
casez ({new_n4452_, new_n5024_})
2'b00 : new_n5943_ = 1'b1;
default : new_n5943_ = 1'b0;
endcase
casez ({new_n2403_, new_n5027_})
2'b11 : new_n5944_ = 1'b1;
default : new_n5944_ = 1'b0;
endcase
casez ({new_n3954_, new_n5063_})
2'b00 : new_n5945_ = 1'b1;
default : new_n5945_ = 1'b0;
endcase
casez ({new_n1777_, new_n5091_})
2'b01 : new_n5946_ = 1'b1;
default : new_n5946_ = 1'b0;
endcase
casez ({new_n3802_, new_n5131_})
2'b00 : new_n5947_ = 1'b1;
default : new_n5947_ = 1'b0;
endcase
casez ({new_n702_, new_n782_})
2'b00 : new_n5948_ = 1'b1;
default : new_n5948_ = 1'b0;
endcase
casez ({new_n3667_, new_n5174_})
2'b10 : new_n5949_ = 1'b1;
default : new_n5949_ = 1'b0;
endcase
casez ({new_n3820_, new_n5194_})
2'b00 : new_n5950_ = 1'b1;
default : new_n5950_ = 1'b0;
endcase
casez ({new_n1763_, new_n5190_})
2'b01 : new_n5951_ = 1'b1;
default : new_n5951_ = 1'b0;
endcase
casez ({new_n1088_, new_n5204_})
2'b01 : new_n5952_ = 1'b1;
default : new_n5952_ = 1'b0;
endcase
casez ({new_n651_, new_n5270_})
2'b01 : new_n5953_ = 1'b1;
default : new_n5953_ = 1'b0;
endcase
casez ({new_n1766_, new_n5295_})
2'b01 : new_n5954_ = 1'b1;
default : new_n5954_ = 1'b0;
endcase
casez ({new_n375_, new_n5296_})
2'b01 : new_n5955_ = 1'b1;
default : new_n5955_ = 1'b0;
endcase
casez ({new_n1250_, new_n5381_})
2'b11 : new_n5956_ = 1'b1;
default : new_n5956_ = 1'b0;
endcase
casez ({new_n4624_, new_n5403_})
2'b00 : new_n5957_ = 1'b1;
default : new_n5957_ = 1'b0;
endcase
casez ({new_n1238_, new_n1990_})
2'b00 : new_n5958_ = 1'b1;
default : new_n5958_ = 1'b0;
endcase
casez ({new_n4972_, new_n5416_})
2'b01 : new_n5959_ = 1'b1;
default : new_n5959_ = 1'b0;
endcase
casez ({new_n2869_, new_n5418_})
2'b01 : new_n5960_ = 1'b1;
default : new_n5960_ = 1'b0;
endcase
casez ({new_n3707_, new_n5427_})
2'b00 : new_n5961_ = 1'b1;
default : new_n5961_ = 1'b0;
endcase
casez ({new_n1237_, new_n1994_})
2'b00 : new_n5962_ = 1'b1;
default : new_n5962_ = 1'b0;
endcase
casez ({new_n3854_, new_n5468_})
2'b01 : new_n5963_ = 1'b1;
default : new_n5963_ = 1'b0;
endcase
casez ({new_n1691_, new_n5479_})
2'b01 : new_n5964_ = 1'b1;
default : new_n5964_ = 1'b0;
endcase
casez ({new_n466_, new_n5486_})
2'b01 : new_n5965_ = 1'b1;
default : new_n5965_ = 1'b0;
endcase
casez ({new_n3060_, new_n5490_})
2'b01 : new_n5966_ = 1'b1;
default : new_n5966_ = 1'b0;
endcase
casez ({new_n2402_, new_n5492_})
2'b11 : new_n5967_ = 1'b1;
default : new_n5967_ = 1'b0;
endcase
casez ({new_n3394_, new_n5500_})
2'b01 : new_n5968_ = 1'b1;
default : new_n5968_ = 1'b0;
endcase
casez ({new_n4275_, new_n5501_})
2'b01 : new_n5969_ = 1'b1;
default : new_n5969_ = 1'b0;
endcase
casez ({new_n1772_, new_n5504_})
2'b01 : new_n5970_ = 1'b1;
default : new_n5970_ = 1'b0;
endcase
casez ({new_n1764_, new_n5523_})
2'b01 : new_n5971_ = 1'b1;
default : new_n5971_ = 1'b0;
endcase
casez ({new_n2312_, new_n5548_})
2'b11 : new_n5972_ = 1'b1;
default : new_n5972_ = 1'b0;
endcase
casez ({new_n4517_, new_n5555_})
2'b01 : new_n5973_ = 1'b1;
default : new_n5973_ = 1'b0;
endcase
casez ({new_n817_, new_n5556_})
2'b01 : new_n5974_ = 1'b1;
default : new_n5974_ = 1'b0;
endcase
casez ({new_n2190_, new_n5574_})
2'b01 : new_n5975_ = 1'b1;
default : new_n5975_ = 1'b0;
endcase
casez ({new_n2168_, new_n5575_})
2'b01 : new_n5976_ = 1'b1;
default : new_n5976_ = 1'b0;
endcase
casez ({new_n2322_, new_n5576_})
2'b01 : new_n5977_ = 1'b1;
default : new_n5977_ = 1'b0;
endcase
casez ({new_n2183_, new_n5577_})
2'b01 : new_n5978_ = 1'b1;
default : new_n5978_ = 1'b0;
endcase
casez ({new_n2225_, new_n5579_})
2'b01 : new_n5979_ = 1'b1;
default : new_n5979_ = 1'b0;
endcase
casez ({new_n474_, new_n5581_})
2'b01 : new_n5980_ = 1'b1;
default : new_n5980_ = 1'b0;
endcase
casez ({new_n2217_, new_n5582_})
2'b01 : new_n5981_ = 1'b1;
default : new_n5981_ = 1'b0;
endcase
casez ({new_n2327_, new_n5585_})
2'b01 : new_n5982_ = 1'b1;
default : new_n5982_ = 1'b0;
endcase
casez ({new_n2258_, new_n5586_})
2'b01 : new_n5983_ = 1'b1;
default : new_n5983_ = 1'b0;
endcase
casez ({new_n1513_, new_n5592_})
2'b11 : new_n5984_ = 1'b1;
default : new_n5984_ = 1'b0;
endcase
casez ({new_n1241_, new_n2041_})
2'b00 : new_n5985_ = 1'b1;
default : new_n5985_ = 1'b0;
endcase
casez ({new_n4489_, new_n5598_})
2'b01 : new_n5986_ = 1'b1;
default : new_n5986_ = 1'b0;
endcase
casez ({new_n4157_, new_n5605_})
2'b01 : new_n5987_ = 1'b1;
default : new_n5987_ = 1'b0;
endcase
casez ({new_n4325_, new_n5608_})
2'b01 : new_n5988_ = 1'b1;
default : new_n5988_ = 1'b0;
endcase
casez ({new_n3866_, new_n5609_})
2'b01 : new_n5989_ = 1'b1;
default : new_n5989_ = 1'b0;
endcase
casez ({new_n4195_, new_n5612_})
2'b01 : new_n5990_ = 1'b1;
default : new_n5990_ = 1'b0;
endcase
casez ({new_n891_, new_n5619_})
2'b01 : new_n5991_ = 1'b1;
default : new_n5991_ = 1'b0;
endcase
casez ({new_n903_, new_n5624_})
2'b01 : new_n5992_ = 1'b1;
default : new_n5992_ = 1'b0;
endcase
casez ({new_n3452_, new_n5629_})
2'b01 : new_n5993_ = 1'b1;
default : new_n5993_ = 1'b0;
endcase
casez ({new_n4681_, new_n5641_})
2'b11 : new_n5994_ = 1'b1;
default : new_n5994_ = 1'b0;
endcase
casez ({new_n5139_, new_n5647_})
2'b01 : new_n5995_ = 1'b1;
default : new_n5995_ = 1'b0;
endcase
casez ({new_n3958_, new_n5651_})
2'b01 : new_n5996_ = 1'b1;
default : new_n5996_ = 1'b0;
endcase
casez ({new_n917_, new_n5652_})
2'b01 : new_n5997_ = 1'b1;
default : new_n5997_ = 1'b0;
endcase
casez ({new_n4781_, new_n5669_})
2'b11 : new_n5998_ = 1'b1;
default : new_n5998_ = 1'b0;
endcase
casez ({new_n3924_, new_n5670_})
2'b01 : new_n5999_ = 1'b1;
default : new_n5999_ = 1'b0;
endcase
casez ({new_n1088_, new_n5671_})
2'b01 : new_n6000_ = 1'b1;
default : new_n6000_ = 1'b0;
endcase
casez ({new_n5472_, new_n5676_})
2'b11 : new_n6001_ = 1'b1;
default : new_n6001_ = 1'b0;
endcase
casez ({new_n3831_, new_n5681_})
2'b01 : new_n6002_ = 1'b1;
default : new_n6002_ = 1'b0;
endcase
casez ({new_n4753_, new_n5686_})
2'b11 : new_n6003_ = 1'b1;
default : new_n6003_ = 1'b0;
endcase
casez ({new_n4067_, new_n5689_})
2'b01 : new_n6004_ = 1'b1;
default : new_n6004_ = 1'b0;
endcase
casez ({new_n2429_, new_n5704_})
2'b01 : new_n6005_ = 1'b1;
default : new_n6005_ = 1'b0;
endcase
casez ({new_n3922_, new_n5715_})
2'b11 : new_n6006_ = 1'b1;
default : new_n6006_ = 1'b0;
endcase
casez ({new_n4773_, new_n5733_})
2'b11 : new_n6007_ = 1'b1;
default : new_n6007_ = 1'b0;
endcase
casez ({new_n1771_, new_n5735_})
2'b01 : new_n6008_ = 1'b1;
default : new_n6008_ = 1'b0;
endcase
casez ({new_n1236_, new_n2052_})
2'b00 : new_n6009_ = 1'b1;
default : new_n6009_ = 1'b0;
endcase
casez ({new_n4847_, new_n5753_})
2'b11 : new_n6010_ = 1'b1;
default : new_n6010_ = 1'b0;
endcase
casez ({new_n5511_, new_n5775_})
2'b11 : new_n6011_ = 1'b1;
default : new_n6011_ = 1'b0;
endcase
casez ({new_n4817_, new_n5805_})
2'b11 : new_n6012_ = 1'b1;
default : new_n6012_ = 1'b0;
endcase
casez ({new_n4828_, new_n5821_})
2'b01 : new_n6013_ = 1'b1;
default : new_n6013_ = 1'b0;
endcase
casez ({new_n5591_, new_n5822_})
2'b11 : new_n6014_ = 1'b1;
default : new_n6014_ = 1'b0;
endcase
casez ({new_n466_, new_n5828_})
2'b01 : new_n6015_ = 1'b1;
default : new_n6015_ = 1'b0;
endcase
casez ({new_n4760_, new_n5832_})
2'b11 : new_n6016_ = 1'b1;
default : new_n6016_ = 1'b0;
endcase
casez ({new_n1830_, new_n5834_})
2'b01 : new_n6017_ = 1'b1;
default : new_n6017_ = 1'b0;
endcase
casez ({new_n4785_, new_n5847_})
2'b11 : new_n6018_ = 1'b1;
default : new_n6018_ = 1'b0;
endcase
casez ({new_n5476_, new_n5855_})
2'b11 : new_n6019_ = 1'b1;
default : new_n6019_ = 1'b0;
endcase
casez ({new_n916_, new_n5865_})
2'b01 : new_n6020_ = 1'b1;
default : new_n6020_ = 1'b0;
endcase
casez ({new_n1086_, new_n5866_})
2'b01 : new_n6021_ = 1'b1;
default : new_n6021_ = 1'b0;
endcase
casez ({new_n1770_, new_n5872_})
2'b01 : new_n6022_ = 1'b1;
default : new_n6022_ = 1'b0;
endcase
casez ({new_n2363_, new_n5874_})
2'b11 : new_n6023_ = 1'b1;
default : new_n6023_ = 1'b0;
endcase
casez ({new_n4965_, new_n5900_})
2'b01 : new_n6024_ = 1'b1;
default : new_n6024_ = 1'b0;
endcase
casez ({new_n2416_, new_n5912_})
2'b11 : new_n6025_ = 1'b1;
default : new_n6025_ = 1'b0;
endcase
casez ({new_n761_, new_n5915_})
2'b11 : new_n6026_ = 1'b1;
default : new_n6026_ = 1'b0;
endcase
casez ({new_n702_, new_n1221_})
2'b00 : new_n6027_ = 1'b1;
default : new_n6027_ = 1'b0;
endcase
casez ({new_n1982_, new_n2175_})
2'b00 : new_n6028_ = 1'b1;
default : new_n6028_ = 1'b0;
endcase
casez ({new_n2065_, new_n2182_})
2'b00 : new_n6029_ = 1'b1;
default : new_n6029_ = 1'b0;
endcase
casez ({new_n2050_, new_n2186_})
2'b00 : new_n6030_ = 1'b1;
default : new_n6030_ = 1'b0;
endcase
casez ({new_n1981_, new_n2195_})
2'b00 : new_n6031_ = 1'b1;
default : new_n6031_ = 1'b0;
endcase
casez ({new_n2185_, new_n2199_})
2'b00 : new_n6032_ = 1'b1;
default : new_n6032_ = 1'b0;
endcase
casez ({new_n1966_, new_n2209_})
2'b00 : new_n6033_ = 1'b1;
default : new_n6033_ = 1'b0;
endcase
casez ({new_n2019_, new_n2210_})
2'b00 : new_n6034_ = 1'b1;
default : new_n6034_ = 1'b0;
endcase
casez ({new_n2032_, new_n2221_})
2'b00 : new_n6035_ = 1'b1;
default : new_n6035_ = 1'b0;
endcase
casez ({new_n2033_, new_n2227_})
2'b00 : new_n6036_ = 1'b1;
default : new_n6036_ = 1'b0;
endcase
casez ({new_n2170_, new_n2228_})
2'b00 : new_n6037_ = 1'b1;
default : new_n6037_ = 1'b0;
endcase
casez ({new_n2086_, new_n2230_})
2'b00 : new_n6038_ = 1'b1;
default : new_n6038_ = 1'b0;
endcase
casez ({new_n1788_, new_n2232_})
2'b00 : new_n6039_ = 1'b1;
default : new_n6039_ = 1'b0;
endcase
casez ({new_n2046_, new_n2234_})
2'b00 : new_n6040_ = 1'b1;
default : new_n6040_ = 1'b0;
endcase
casez ({new_n2057_, new_n2235_})
2'b00 : new_n6041_ = 1'b1;
default : new_n6041_ = 1'b0;
endcase
casez ({new_n2233_, new_n2236_})
2'b00 : new_n6042_ = 1'b1;
default : new_n6042_ = 1'b0;
endcase
casez ({new_n2176_, new_n2250_})
2'b00 : new_n6043_ = 1'b1;
default : new_n6043_ = 1'b0;
endcase
casez ({new_n1971_, new_n2251_})
2'b00 : new_n6044_ = 1'b1;
default : new_n6044_ = 1'b0;
endcase
casez ({new_n2238_, new_n2253_})
2'b00 : new_n6045_ = 1'b1;
default : new_n6045_ = 1'b0;
endcase
casez ({new_n2248_, new_n2255_})
2'b00 : new_n6046_ = 1'b1;
default : new_n6046_ = 1'b0;
endcase
casez ({new_n2247_, new_n2272_})
2'b00 : new_n6047_ = 1'b1;
default : new_n6047_ = 1'b0;
endcase
casez ({new_n2207_, new_n2276_})
2'b00 : new_n6048_ = 1'b1;
default : new_n6048_ = 1'b0;
endcase
casez ({new_n1988_, new_n2288_})
2'b00 : new_n6049_ = 1'b1;
default : new_n6049_ = 1'b0;
endcase
casez ({new_n2198_, new_n2291_})
2'b00 : new_n6050_ = 1'b1;
default : new_n6050_ = 1'b0;
endcase
casez ({new_n914_, new_n1322_})
2'b00 : new_n6051_ = 1'b1;
default : new_n6051_ = 1'b0;
endcase
casez ({new_n2283_, new_n2300_})
2'b00 : new_n6052_ = 1'b1;
default : new_n6052_ = 1'b0;
endcase
casez ({new_n2184_, new_n2303_})
2'b00 : new_n6053_ = 1'b1;
default : new_n6053_ = 1'b0;
endcase
casez ({new_n2053_, new_n2307_})
2'b00 : new_n6054_ = 1'b1;
default : new_n6054_ = 1'b0;
endcase
casez ({new_n2093_, new_n2320_})
2'b00 : new_n6055_ = 1'b1;
default : new_n6055_ = 1'b0;
endcase
casez ({new_n2262_, new_n2323_})
2'b00 : new_n6056_ = 1'b1;
default : new_n6056_ = 1'b0;
endcase
casez ({new_n2089_, new_n2330_})
2'b00 : new_n6057_ = 1'b1;
default : new_n6057_ = 1'b0;
endcase
casez ({new_n2271_, new_n2331_})
2'b00 : new_n6058_ = 1'b1;
default : new_n6058_ = 1'b0;
endcase
casez ({new_n2281_, new_n2333_})
2'b00 : new_n6059_ = 1'b1;
default : new_n6059_ = 1'b0;
endcase
casez ({new_n1145_, new_n2338_})
2'b01 : new_n6060_ = 1'b1;
default : new_n6060_ = 1'b0;
endcase
casez ({new_n596_, new_n880_})
2'b00 : new_n6061_ = 1'b1;
default : new_n6061_ = 1'b0;
endcase
casez ({new_n1384_, new_n2402_})
2'b01 : new_n6062_ = 1'b1;
default : new_n6062_ = 1'b0;
endcase
casez ({new_n1858_, new_n2403_})
2'b01 : new_n6063_ = 1'b1;
default : new_n6063_ = 1'b0;
endcase
casez ({new_n1519_, new_n2408_})
2'b01 : new_n6064_ = 1'b1;
default : new_n6064_ = 1'b0;
endcase
casez ({new_n871_, new_n2425_})
2'b01 : new_n6065_ = 1'b1;
default : new_n6065_ = 1'b0;
endcase
casez ({new_n644_, new_n2426_})
2'b01 : new_n6066_ = 1'b1;
default : new_n6066_ = 1'b0;
endcase
casez ({new_n1615_, new_n2426_})
2'b01 : new_n6067_ = 1'b1;
default : new_n6067_ = 1'b0;
endcase
casez ({new_n521_, new_n914_})
2'b00 : new_n6068_ = 1'b1;
default : new_n6068_ = 1'b0;
endcase
casez ({new_n1085_, new_n2558_})
2'b00 : new_n6069_ = 1'b1;
default : new_n6069_ = 1'b0;
endcase
casez ({new_n1787_, new_n2581_})
2'b00 : new_n6070_ = 1'b1;
default : new_n6070_ = 1'b0;
endcase
casez ({new_n1088_, new_n2604_})
2'b00 : new_n6071_ = 1'b1;
default : new_n6071_ = 1'b0;
endcase
casez ({new_n596_, new_n2610_})
2'b00 : new_n6072_ = 1'b1;
default : new_n6072_ = 1'b0;
endcase
casez ({new_n1078_, new_n2653_})
2'b00 : new_n6073_ = 1'b1;
default : new_n6073_ = 1'b0;
endcase
casez ({new_n375_, new_n945_})
2'b00 : new_n6074_ = 1'b1;
default : new_n6074_ = 1'b0;
endcase
casez ({new_n1528_, new_n2671_})
2'b10 : new_n6075_ = 1'b1;
default : new_n6075_ = 1'b0;
endcase
casez ({new_n1519_, new_n2731_})
2'b00 : new_n6076_ = 1'b1;
default : new_n6076_ = 1'b0;
endcase
casez ({new_n595_, new_n2740_})
2'b00 : new_n6077_ = 1'b1;
default : new_n6077_ = 1'b0;
endcase
casez ({new_n762_, new_n1490_})
2'b00 : new_n6078_ = 1'b1;
default : new_n6078_ = 1'b0;
endcase
casez ({new_n1079_, new_n1500_})
2'b00 : new_n6079_ = 1'b1;
default : new_n6079_ = 1'b0;
endcase
casez ({new_n1510_, new_n2820_})
2'b00 : new_n6080_ = 1'b1;
default : new_n6080_ = 1'b0;
endcase
casez ({new_n1080_, new_n2823_})
2'b00 : new_n6081_ = 1'b1;
default : new_n6081_ = 1'b0;
endcase
casez ({new_n1199_, new_n1508_})
2'b00 : new_n6082_ = 1'b1;
default : new_n6082_ = 1'b0;
endcase
casez ({new_n610_, new_n1522_})
2'b00 : new_n6083_ = 1'b1;
default : new_n6083_ = 1'b0;
endcase
casez ({new_n566_, new_n1528_})
2'b01 : new_n6084_ = 1'b1;
default : new_n6084_ = 1'b0;
endcase
casez ({new_n577_, new_n651_})
2'b00 : new_n6085_ = 1'b1;
default : new_n6085_ = 1'b0;
endcase
casez ({new_n1517_, new_n1562_})
2'b00 : new_n6086_ = 1'b1;
default : new_n6086_ = 1'b0;
endcase
casez ({new_n375_, new_n2958_})
2'b00 : new_n6087_ = 1'b1;
default : new_n6087_ = 1'b0;
endcase
casez ({new_n1766_, new_n3312_})
2'b00 : new_n6088_ = 1'b1;
default : new_n6088_ = 1'b0;
endcase
casez ({new_n374_, new_n1037_})
2'b00 : new_n6089_ = 1'b1;
default : new_n6089_ = 1'b0;
endcase
casez ({new_n464_, new_n700_})
2'b00 : new_n6090_ = 1'b1;
default : new_n6090_ = 1'b0;
endcase
casez ({new_n1771_, new_n3648_})
2'b01 : new_n6091_ = 1'b1;
default : new_n6091_ = 1'b0;
endcase
casez ({new_n1536_, new_n3709_})
2'b11 : new_n6092_ = 1'b1;
default : new_n6092_ = 1'b0;
endcase
casez ({new_n1763_, new_n3814_})
2'b00 : new_n6093_ = 1'b1;
default : new_n6093_ = 1'b0;
endcase
casez ({new_n1517_, new_n3883_})
2'b01 : new_n6094_ = 1'b1;
default : new_n6094_ = 1'b0;
endcase
casez ({new_n1507_, new_n3896_})
2'b00 : new_n6095_ = 1'b1;
default : new_n6095_ = 1'b0;
endcase
casez ({new_n807_, new_n1075_})
2'b00 : new_n6096_ = 1'b1;
default : new_n6096_ = 1'b0;
endcase
casez ({new_n702_, new_n3996_})
2'b00 : new_n6097_ = 1'b1;
default : new_n6097_ = 1'b0;
endcase
casez ({new_n843_, new_n1080_})
2'b00 : new_n6098_ = 1'b1;
default : new_n6098_ = 1'b0;
endcase
casez ({new_n521_, new_n1081_})
2'b00 : new_n6099_ = 1'b1;
default : new_n6099_ = 1'b0;
endcase
casez ({new_n817_, new_n4026_})
2'b00 : new_n6100_ = 1'b1;
default : new_n6100_ = 1'b0;
endcase
casez ({new_n778_, new_n1083_})
2'b00 : new_n6101_ = 1'b1;
default : new_n6101_ = 1'b0;
endcase
casez ({new_n331_, new_n4065_})
2'b01 : new_n6102_ = 1'b1;
default : new_n6102_ = 1'b0;
endcase
casez ({new_n1629_, new_n1773_})
2'b00 : new_n6103_ = 1'b1;
default : new_n6103_ = 1'b0;
endcase
casez ({new_n2869_, new_n4098_})
2'b01 : new_n6104_ = 1'b1;
default : new_n6104_ = 1'b0;
endcase
casez ({new_n798_, new_n1777_})
2'b00 : new_n6105_ = 1'b1;
default : new_n6105_ = 1'b0;
endcase
casez ({new_n914_, new_n4137_})
2'b01 : new_n6106_ = 1'b1;
default : new_n6106_ = 1'b0;
endcase
casez ({new_n1571_, new_n1787_})
2'b00 : new_n6107_ = 1'b1;
default : new_n6107_ = 1'b0;
endcase
casez ({new_n1611_, new_n1787_})
2'b00 : new_n6108_ = 1'b1;
default : new_n6108_ = 1'b0;
endcase
casez ({new_n626_, new_n4245_})
2'b01 : new_n6109_ = 1'b1;
default : new_n6109_ = 1'b0;
endcase
casez ({new_n2408_, new_n4290_})
2'b11 : new_n6110_ = 1'b1;
default : new_n6110_ = 1'b0;
endcase
casez ({new_n762_, new_n4379_})
2'b01 : new_n6111_ = 1'b1;
default : new_n6111_ = 1'b0;
endcase
casez ({new_n1787_, new_n4408_})
2'b01 : new_n6112_ = 1'b1;
default : new_n6112_ = 1'b0;
endcase
casez ({new_n1510_, new_n1844_})
2'b00 : new_n6113_ = 1'b1;
default : new_n6113_ = 1'b0;
endcase
casez ({new_n762_, new_n4544_})
2'b01 : new_n6114_ = 1'b1;
default : new_n6114_ = 1'b0;
endcase
casez ({new_n1776_, new_n1860_})
2'b00 : new_n6115_ = 1'b1;
default : new_n6115_ = 1'b0;
endcase
casez ({new_n817_, new_n1865_})
2'b00 : new_n6116_ = 1'b1;
default : new_n6116_ = 1'b0;
endcase
casez ({new_n686_, new_n4672_})
2'b00 : new_n6117_ = 1'b1;
default : new_n6117_ = 1'b0;
endcase
casez ({new_n1761_, new_n4757_})
2'b01 : new_n6118_ = 1'b1;
default : new_n6118_ = 1'b0;
endcase
casez ({new_n1507_, new_n4765_})
2'b01 : new_n6119_ = 1'b1;
default : new_n6119_ = 1'b0;
endcase
casez ({new_n2845_, new_n4775_})
2'b00 : new_n6120_ = 1'b1;
default : new_n6120_ = 1'b0;
endcase
casez ({new_n596_, new_n4814_})
2'b01 : new_n6121_ = 1'b1;
default : new_n6121_ = 1'b0;
endcase
casez ({new_n468_, new_n4841_})
2'b00 : new_n6122_ = 1'b1;
default : new_n6122_ = 1'b0;
endcase
casez ({new_n287_, new_n420_, new_n5043_})
3'b11? : new_n6123_ = 1'b1;
3'b??1 : new_n6123_ = 1'b1;
default : new_n6123_ = 1'b0;
endcase
casez ({new_n375_, new_n476_, new_n2820_})
3'b11? : new_n6124_ = 1'b1;
3'b??1 : new_n6124_ = 1'b1;
default : new_n6124_ = 1'b0;
endcase
casez ({x[1], new_n375_, new_n1072_})
3'b01? : new_n6125_ = 1'b1;
3'b??1 : new_n6125_ = 1'b1;
default : new_n6125_ = 1'b0;
endcase
casez ({new_n252_, new_n749_, new_n1844_})
3'b01? : new_n6126_ = 1'b1;
3'b??1 : new_n6126_ = 1'b1;
default : new_n6126_ = 1'b0;
endcase
casez ({new_n327_, new_n467_})
2'b00 : new_n6127_ = 1'b1;
default : new_n6127_ = 1'b0;
endcase
casez ({new_n85_, new_n374_})
2'b11 : new_n6128_ = 1'b1;
default : new_n6128_ = 1'b0;
endcase
casez ({new_n224_, new_n1529_})
2'b10 : new_n6129_ = 1'b1;
default : new_n6129_ = 1'b0;
endcase
casez ({new_n85_, new_n761_})
2'b10 : new_n6130_ = 1'b1;
default : new_n6130_ = 1'b0;
endcase
casez ({new_n1254_, new_n1903_})
2'b00 : new_n6131_ = 1'b1;
default : new_n6131_ = 1'b0;
endcase
casez ({new_n614_, new_n5145_})
2'b01 : new_n6132_ = 1'b1;
default : new_n6132_ = 1'b0;
endcase
casez ({new_n1249_, new_n1984_})
2'b00 : new_n6133_ = 1'b1;
default : new_n6133_ = 1'b0;
endcase
casez ({new_n1254_, new_n5419_})
2'b01 : new_n6134_ = 1'b1;
default : new_n6134_ = 1'b0;
endcase
casez ({new_n1242_, new_n5580_})
2'b00 : new_n6135_ = 1'b1;
default : new_n6135_ = 1'b0;
endcase
casez ({new_n4075_, new_n5778_})
2'b00 : new_n6136_ = 1'b1;
default : new_n6136_ = 1'b0;
endcase
casez ({new_n1089_, new_n5863_})
2'b01 : new_n6137_ = 1'b1;
default : new_n6137_ = 1'b0;
endcase
casez ({new_n1785_, new_n5882_})
2'b01 : new_n6138_ = 1'b1;
default : new_n6138_ = 1'b0;
endcase
casez ({new_n761_, new_n5937_})
2'b11 : new_n6139_ = 1'b1;
default : new_n6139_ = 1'b0;
endcase
casez ({new_n2852_, new_n5975_})
2'b01 : new_n6140_ = 1'b1;
default : new_n6140_ = 1'b0;
endcase
casez ({new_n2390_, new_n5977_})
2'b01 : new_n6141_ = 1'b1;
default : new_n6141_ = 1'b0;
endcase
casez ({new_n2401_, new_n5978_})
2'b01 : new_n6142_ = 1'b1;
default : new_n6142_ = 1'b0;
endcase
casez ({new_n2419_, new_n5979_})
2'b01 : new_n6143_ = 1'b1;
default : new_n6143_ = 1'b0;
endcase
casez ({new_n2397_, new_n5981_})
2'b01 : new_n6144_ = 1'b1;
default : new_n6144_ = 1'b0;
endcase
casez ({new_n2396_, new_n5983_})
2'b01 : new_n6145_ = 1'b1;
default : new_n6145_ = 1'b0;
endcase
casez ({new_n2428_, new_n5985_})
2'b01 : new_n6146_ = 1'b1;
default : new_n6146_ = 1'b0;
endcase
casez ({new_n1780_, new_n5989_})
2'b01 : new_n6147_ = 1'b1;
default : new_n6147_ = 1'b0;
endcase
casez ({new_n2863_, new_n6009_})
2'b01 : new_n6148_ = 1'b1;
default : new_n6148_ = 1'b0;
endcase
casez ({new_n1533_, new_n6016_})
2'b11 : new_n6149_ = 1'b1;
default : new_n6149_ = 1'b0;
endcase
casez ({new_n2386_, new_n6028_})
2'b01 : new_n6150_ = 1'b1;
default : new_n6150_ = 1'b0;
endcase
casez ({new_n2854_, new_n6029_})
2'b01 : new_n6151_ = 1'b1;
default : new_n6151_ = 1'b0;
endcase
casez ({new_n2286_, new_n6034_})
2'b01 : new_n6152_ = 1'b1;
default : new_n6152_ = 1'b0;
endcase
casez ({new_n2423_, new_n6035_})
2'b01 : new_n6153_ = 1'b1;
default : new_n6153_ = 1'b0;
endcase
casez ({new_n2266_, new_n6036_})
2'b01 : new_n6154_ = 1'b1;
default : new_n6154_ = 1'b0;
endcase
casez ({new_n2345_, new_n6037_})
2'b01 : new_n6155_ = 1'b1;
default : new_n6155_ = 1'b0;
endcase
casez ({new_n2405_, new_n6038_})
2'b01 : new_n6156_ = 1'b1;
default : new_n6156_ = 1'b0;
endcase
casez ({new_n2415_, new_n6039_})
2'b01 : new_n6157_ = 1'b1;
default : new_n6157_ = 1'b0;
endcase
casez ({new_n5976_, new_n6040_})
2'b11 : new_n6158_ = 1'b1;
default : new_n6158_ = 1'b0;
endcase
casez ({new_n2348_, new_n6041_})
2'b01 : new_n6159_ = 1'b1;
default : new_n6159_ = 1'b0;
endcase
casez ({new_n2349_, new_n6042_})
2'b01 : new_n6160_ = 1'b1;
default : new_n6160_ = 1'b0;
endcase
casez ({new_n2392_, new_n6043_})
2'b01 : new_n6161_ = 1'b1;
default : new_n6161_ = 1'b0;
endcase
casez ({new_n2861_, new_n6047_})
2'b01 : new_n6162_ = 1'b1;
default : new_n6162_ = 1'b0;
endcase
casez ({new_n2355_, new_n6050_})
2'b01 : new_n6163_ = 1'b1;
default : new_n6163_ = 1'b0;
endcase
casez ({new_n594_, new_n6051_})
2'b01 : new_n6164_ = 1'b1;
default : new_n6164_ = 1'b0;
endcase
casez ({new_n6045_, new_n6052_})
2'b11 : new_n6165_ = 1'b1;
default : new_n6165_ = 1'b0;
endcase
casez ({new_n2347_, new_n6054_})
2'b01 : new_n6166_ = 1'b1;
default : new_n6166_ = 1'b0;
endcase
casez ({new_n705_, new_n850_})
2'b00 : new_n6167_ = 1'b1;
default : new_n6167_ = 1'b0;
endcase
casez ({new_n6046_, new_n6058_})
2'b11 : new_n6168_ = 1'b1;
default : new_n6168_ = 1'b0;
endcase
casez ({new_n4268_, new_n6064_})
2'b01 : new_n6169_ = 1'b1;
default : new_n6169_ = 1'b0;
endcase
casez ({new_n4840_, new_n6071_})
2'b01 : new_n6170_ = 1'b1;
default : new_n6170_ = 1'b0;
endcase
casez ({new_n1778_, new_n2224_})
2'b01 : new_n6171_ = 1'b1;
default : new_n6171_ = 1'b0;
endcase
casez ({new_n1247_, new_n2316_})
2'b00 : new_n6172_ = 1'b1;
default : new_n6172_ = 1'b0;
endcase
casez ({new_n2060_, new_n2340_})
2'b00 : new_n6173_ = 1'b1;
default : new_n6173_ = 1'b0;
endcase
casez ({new_n2205_, new_n2342_})
2'b00 : new_n6174_ = 1'b1;
default : new_n6174_ = 1'b0;
endcase
casez ({new_n1781_, new_n2343_})
2'b00 : new_n6175_ = 1'b1;
default : new_n6175_ = 1'b0;
endcase
casez ({new_n2284_, new_n2344_})
2'b00 : new_n6176_ = 1'b1;
default : new_n6176_ = 1'b0;
endcase
casez ({new_n2202_, new_n2346_})
2'b00 : new_n6177_ = 1'b1;
default : new_n6177_ = 1'b0;
endcase
casez ({new_n2213_, new_n2351_})
2'b00 : new_n6178_ = 1'b1;
default : new_n6178_ = 1'b0;
endcase
casez ({new_n2315_, new_n2352_})
2'b00 : new_n6179_ = 1'b1;
default : new_n6179_ = 1'b0;
endcase
casez ({new_n2325_, new_n2354_})
2'b00 : new_n6180_ = 1'b1;
default : new_n6180_ = 1'b0;
endcase
casez ({new_n2274_, new_n2356_})
2'b00 : new_n6181_ = 1'b1;
default : new_n6181_ = 1'b0;
endcase
casez ({new_n2306_, new_n2357_})
2'b00 : new_n6182_ = 1'b1;
default : new_n6182_ = 1'b0;
endcase
casez ({new_n2191_, new_n2364_})
2'b00 : new_n6183_ = 1'b1;
default : new_n6183_ = 1'b0;
endcase
casez ({new_n2043_, new_n2376_})
2'b00 : new_n6184_ = 1'b1;
default : new_n6184_ = 1'b0;
endcase
casez ({new_n2054_, new_n2383_})
2'b00 : new_n6185_ = 1'b1;
default : new_n6185_ = 1'b0;
endcase
casez ({new_n731_, new_n2385_})
2'b00 : new_n6186_ = 1'b1;
default : new_n6186_ = 1'b0;
endcase
casez ({new_n2285_, new_n2410_})
2'b00 : new_n6187_ = 1'b1;
default : new_n6187_ = 1'b0;
endcase
casez ({new_n2167_, new_n2411_})
2'b00 : new_n6188_ = 1'b1;
default : new_n6188_ = 1'b0;
endcase
casez ({new_n2077_, new_n2417_})
2'b00 : new_n6189_ = 1'b1;
default : new_n6189_ = 1'b0;
endcase
casez ({new_n2377_, new_n2427_})
2'b00 : new_n6190_ = 1'b1;
default : new_n6190_ = 1'b0;
endcase
casez ({new_n819_, new_n2473_})
2'b01 : new_n6191_ = 1'b1;
default : new_n6191_ = 1'b0;
endcase
casez ({new_n384_, new_n614_})
2'b00 : new_n6192_ = 1'b1;
default : new_n6192_ = 1'b0;
endcase
casez ({new_n614_, new_n2593_})
2'b00 : new_n6193_ = 1'b1;
default : new_n6193_ = 1'b0;
endcase
casez ({new_n1254_, new_n2614_})
2'b00 : new_n6194_ = 1'b1;
default : new_n6194_ = 1'b0;
endcase
casez ({new_n2087_, new_n2856_})
2'b00 : new_n6195_ = 1'b1;
default : new_n6195_ = 1'b0;
endcase
casez ({new_n2361_, new_n2865_})
2'b00 : new_n6196_ = 1'b1;
default : new_n6196_ = 1'b0;
endcase
casez ({new_n2422_, new_n2871_})
2'b01 : new_n6197_ = 1'b1;
default : new_n6197_ = 1'b0;
endcase
casez ({new_n614_, new_n1014_})
2'b00 : new_n6198_ = 1'b1;
default : new_n6198_ = 1'b0;
endcase
casez ({new_n1341_, new_n1778_})
2'b00 : new_n6199_ = 1'b1;
default : new_n6199_ = 1'b0;
endcase
casez ({new_n510_, new_n1782_})
2'b00 : new_n6200_ = 1'b1;
default : new_n6200_ = 1'b0;
endcase
casez ({new_n837_, new_n1785_})
2'b00 : new_n6201_ = 1'b1;
default : new_n6201_ = 1'b0;
endcase
casez ({new_n1783_, new_n4347_})
2'b01 : new_n6202_ = 1'b1;
default : new_n6202_ = 1'b0;
endcase
casez ({new_n1782_, new_n1845_})
2'b00 : new_n6203_ = 1'b1;
default : new_n6203_ = 1'b0;
endcase
casez ({new_n614_, new_n1121_})
2'b00 : new_n6204_ = 1'b1;
default : new_n6204_ = 1'b0;
endcase
casez ({new_n275_, new_n1541_, new_n1780_})
3'b10? : new_n6205_ = 1'b1;
3'b??1 : new_n6205_ = 1'b1;
default : new_n6205_ = 1'b0;
endcase
casez ({new_n1790_, new_n5939_})
2'b01 : new_n6206_ = 1'b1;
default : new_n6206_ = 1'b0;
endcase
casez ({new_n1253_, new_n2097_})
2'b00 : new_n6207_ = 1'b1;
default : new_n6207_ = 1'b0;
endcase
casez ({new_n2466_, new_n5982_})
2'b01 : new_n6208_ = 1'b1;
default : new_n6208_ = 1'b0;
endcase
casez ({new_n2889_, new_n6048_})
2'b11 : new_n6209_ = 1'b1;
default : new_n6209_ = 1'b0;
endcase
casez ({new_n2432_, new_n6056_})
2'b01 : new_n6210_ = 1'b1;
default : new_n6210_ = 1'b0;
endcase
casez ({new_n6030_, new_n6140_})
2'b11 : new_n6211_ = 1'b1;
default : new_n6211_ = 1'b0;
endcase
casez ({new_n2458_, new_n6141_})
2'b01 : new_n6212_ = 1'b1;
default : new_n6212_ = 1'b0;
endcase
casez ({new_n2463_, new_n6142_})
2'b01 : new_n6213_ = 1'b1;
default : new_n6213_ = 1'b0;
endcase
casez ({new_n2460_, new_n6143_})
2'b01 : new_n6214_ = 1'b1;
default : new_n6214_ = 1'b0;
endcase
casez ({new_n2469_, new_n6144_})
2'b01 : new_n6215_ = 1'b1;
default : new_n6215_ = 1'b0;
endcase
casez ({new_n2256_, new_n6146_})
2'b01 : new_n6216_ = 1'b1;
default : new_n6216_ = 1'b0;
endcase
casez ({new_n6059_, new_n6151_})
2'b11 : new_n6217_ = 1'b1;
default : new_n6217_ = 1'b0;
endcase
casez ({new_n2462_, new_n6154_})
2'b01 : new_n6218_ = 1'b1;
default : new_n6218_ = 1'b0;
endcase
casez ({new_n2890_, new_n6155_})
2'b11 : new_n6219_ = 1'b1;
default : new_n6219_ = 1'b0;
endcase
casez ({new_n2295_, new_n6156_})
2'b01 : new_n6220_ = 1'b1;
default : new_n6220_ = 1'b0;
endcase
casez ({new_n2280_, new_n6157_})
2'b01 : new_n6221_ = 1'b1;
default : new_n6221_ = 1'b0;
endcase
casez ({new_n2470_, new_n6158_})
2'b01 : new_n6222_ = 1'b1;
default : new_n6222_ = 1'b0;
endcase
casez ({new_n2471_, new_n6159_})
2'b01 : new_n6223_ = 1'b1;
default : new_n6223_ = 1'b0;
endcase
casez ({new_n2459_, new_n6160_})
2'b01 : new_n6224_ = 1'b1;
default : new_n6224_ = 1'b0;
endcase
casez ({new_n2464_, new_n6161_})
2'b01 : new_n6225_ = 1'b1;
default : new_n6225_ = 1'b0;
endcase
casez ({new_n2389_, new_n6163_})
2'b01 : new_n6226_ = 1'b1;
default : new_n6226_ = 1'b0;
endcase
casez ({new_n2375_, new_n6166_})
2'b01 : new_n6227_ = 1'b1;
default : new_n6227_ = 1'b0;
endcase
casez ({new_n2413_, new_n6173_})
2'b01 : new_n6228_ = 1'b1;
default : new_n6228_ = 1'b0;
endcase
casez ({new_n2882_, new_n6176_})
2'b01 : new_n6229_ = 1'b1;
default : new_n6229_ = 1'b0;
endcase
casez ({new_n2864_, new_n6177_})
2'b01 : new_n6230_ = 1'b1;
default : new_n6230_ = 1'b0;
endcase
casez ({new_n2862_, new_n6178_})
2'b01 : new_n6231_ = 1'b1;
default : new_n6231_ = 1'b0;
endcase
casez ({new_n2866_, new_n6179_})
2'b01 : new_n6232_ = 1'b1;
default : new_n6232_ = 1'b0;
endcase
casez ({new_n2868_, new_n6180_})
2'b01 : new_n6233_ = 1'b1;
default : new_n6233_ = 1'b0;
endcase
casez ({new_n2373_, new_n6181_})
2'b01 : new_n6234_ = 1'b1;
default : new_n6234_ = 1'b0;
endcase
casez ({new_n2414_, new_n6183_})
2'b01 : new_n6235_ = 1'b1;
default : new_n6235_ = 1'b0;
endcase
casez ({new_n6133_, new_n6186_})
2'b11 : new_n6236_ = 1'b1;
default : new_n6236_ = 1'b0;
endcase
casez ({new_n2857_, new_n6189_})
2'b01 : new_n6237_ = 1'b1;
default : new_n6237_ = 1'b0;
endcase
casez ({new_n2468_, new_n6190_})
2'b01 : new_n6238_ = 1'b1;
default : new_n6238_ = 1'b0;
endcase
casez ({new_n6172_, new_n6196_})
2'b11 : new_n6239_ = 1'b1;
default : new_n6239_ = 1'b0;
endcase
casez ({new_n6182_, new_n6197_})
2'b11 : new_n6240_ = 1'b1;
default : new_n6240_ = 1'b0;
endcase
casez ({new_n2393_, new_n2435_})
2'b00 : new_n6241_ = 1'b1;
default : new_n6241_ = 1'b0;
endcase
casez ({new_n2433_, new_n2436_})
2'b00 : new_n6242_ = 1'b1;
default : new_n6242_ = 1'b0;
endcase
casez ({new_n2371_, new_n2446_})
2'b00 : new_n6243_ = 1'b1;
default : new_n6243_ = 1'b0;
endcase
casez ({new_n2404_, new_n2447_})
2'b00 : new_n6244_ = 1'b1;
default : new_n6244_ = 1'b0;
endcase
casez ({new_n2443_, new_n2448_})
2'b00 : new_n6245_ = 1'b1;
default : new_n6245_ = 1'b0;
endcase
casez ({new_n2388_, new_n2451_})
2'b00 : new_n6246_ = 1'b1;
default : new_n6246_ = 1'b0;
endcase
casez ({new_n2378_, new_n2453_})
2'b00 : new_n6247_ = 1'b1;
default : new_n6247_ = 1'b0;
endcase
casez ({new_n2421_, new_n2457_})
2'b00 : new_n6248_ = 1'b1;
default : new_n6248_ = 1'b0;
endcase
casez ({new_n2454_, new_n2474_})
2'b00 : new_n6249_ = 1'b1;
default : new_n6249_ = 1'b0;
endcase
casez ({new_n2214_, new_n2873_})
2'b00 : new_n6250_ = 1'b1;
default : new_n6250_ = 1'b0;
endcase
casez ({new_n2212_, new_n2874_})
2'b00 : new_n6251_ = 1'b1;
default : new_n6251_ = 1'b0;
endcase
casez ({new_n2201_, new_n2875_})
2'b00 : new_n6252_ = 1'b1;
default : new_n6252_ = 1'b0;
endcase
casez ({new_n2412_, new_n2876_})
2'b00 : new_n6253_ = 1'b1;
default : new_n6253_ = 1'b0;
endcase
casez ({new_n2400_, new_n2878_})
2'b00 : new_n6254_ = 1'b1;
default : new_n6254_ = 1'b0;
endcase
casez ({new_n2321_, new_n2879_})
2'b00 : new_n6255_ = 1'b1;
default : new_n6255_ = 1'b0;
endcase
casez ({new_n2269_, new_n2881_})
2'b00 : new_n6256_ = 1'b1;
default : new_n6256_ = 1'b0;
endcase
casez ({new_n2372_, new_n2886_})
2'b00 : new_n6257_ = 1'b1;
default : new_n6257_ = 1'b0;
endcase
casez ({new_n1793_, new_n6053_})
2'b01 : new_n6258_ = 1'b1;
default : new_n6258_ = 1'b0;
endcase
casez ({new_n2484_, new_n6145_})
2'b01 : new_n6259_ = 1'b1;
default : new_n6259_ = 1'b0;
endcase
casez ({new_n2891_, new_n6168_})
2'b01 : new_n6260_ = 1'b1;
default : new_n6260_ = 1'b0;
endcase
casez ({new_n6148_, new_n6209_})
2'b11 : new_n6261_ = 1'b1;
default : new_n6261_ = 1'b0;
endcase
casez ({new_n2486_, new_n6212_})
2'b01 : new_n6262_ = 1'b1;
default : new_n6262_ = 1'b0;
endcase
casez ({new_n6165_, new_n6213_})
2'b11 : new_n6263_ = 1'b1;
default : new_n6263_ = 1'b0;
endcase
casez ({new_n2240_, new_n6214_})
2'b01 : new_n6264_ = 1'b1;
default : new_n6264_ = 1'b0;
endcase
casez ({new_n6175_, new_n6218_})
2'b11 : new_n6265_ = 1'b1;
default : new_n6265_ = 1'b0;
endcase
casez ({new_n6219_, new_n6224_})
2'b11 : new_n6266_ = 1'b1;
default : new_n6266_ = 1'b0;
endcase
casez ({new_n6215_, new_n6226_})
2'b11 : new_n6267_ = 1'b1;
default : new_n6267_ = 1'b0;
endcase
casez ({new_n2487_, new_n6227_})
2'b01 : new_n6268_ = 1'b1;
default : new_n6268_ = 1'b0;
endcase
casez ({new_n2366_, new_n6229_})
2'b01 : new_n6269_ = 1'b1;
default : new_n6269_ = 1'b0;
endcase
casez ({new_n2887_, new_n6241_})
2'b01 : new_n6270_ = 1'b1;
default : new_n6270_ = 1'b0;
endcase
casez ({new_n2475_, new_n6243_})
2'b01 : new_n6271_ = 1'b1;
default : new_n6271_ = 1'b0;
endcase
casez ({new_n2481_, new_n6244_})
2'b01 : new_n6272_ = 1'b1;
default : new_n6272_ = 1'b0;
endcase
casez ({new_n2450_, new_n6245_})
2'b01 : new_n6273_ = 1'b1;
default : new_n6273_ = 1'b0;
endcase
casez ({new_n2898_, new_n6247_})
2'b01 : new_n6274_ = 1'b1;
default : new_n6274_ = 1'b0;
endcase
casez ({new_n2480_, new_n6249_})
2'b01 : new_n6275_ = 1'b1;
default : new_n6275_ = 1'b0;
endcase
casez ({new_n2467_, new_n2477_})
2'b00 : new_n6276_ = 1'b1;
default : new_n6276_ = 1'b0;
endcase
casez ({new_n2438_, new_n2478_})
2'b00 : new_n6277_ = 1'b1;
default : new_n6277_ = 1'b0;
endcase
casez ({new_n2485_, new_n2489_})
2'b00 : new_n6278_ = 1'b1;
default : new_n6278_ = 1'b0;
endcase
casez ({new_n2252_, new_n2490_})
2'b00 : new_n6279_ = 1'b1;
default : new_n6279_ = 1'b0;
endcase
casez ({new_n2360_, new_n2892_})
2'b00 : new_n6280_ = 1'b1;
default : new_n6280_ = 1'b0;
endcase
casez ({new_n2449_, new_n2893_})
2'b00 : new_n6281_ = 1'b1;
default : new_n6281_ = 1'b0;
endcase
casez ({new_n2445_, new_n2897_})
2'b00 : new_n6282_ = 1'b1;
default : new_n6282_ = 1'b0;
endcase
casez ({new_n1794_, new_n6057_})
2'b01 : new_n6283_ = 1'b1;
default : new_n6283_ = 1'b0;
endcase
casez ({new_n922_, new_n6207_})
2'b01 : new_n6284_ = 1'b1;
default : new_n6284_ = 1'b0;
endcase
casez ({new_n2492_, new_n6223_})
2'b01 : new_n6285_ = 1'b1;
default : new_n6285_ = 1'b0;
endcase
casez ({new_n2902_, new_n6242_})
2'b01 : new_n6286_ = 1'b1;
default : new_n6286_ = 1'b0;
endcase
casez ({new_n6222_, new_n6260_})
2'b11 : new_n6287_ = 1'b1;
default : new_n6287_ = 1'b0;
endcase
casez ({new_n6262_, new_n6264_})
2'b11 : new_n6288_ = 1'b1;
default : new_n6288_ = 1'b0;
endcase
casez ({new_n6263_, new_n6266_})
2'b11 : new_n6289_ = 1'b1;
default : new_n6289_ = 1'b0;
endcase
casez ({new_n2894_, new_n6273_})
2'b01 : new_n6290_ = 1'b1;
default : new_n6290_ = 1'b0;
endcase
casez ({new_n6275_, new_n6278_})
2'b11 : new_n6291_ = 1'b1;
default : new_n6291_ = 1'b0;
endcase
casez ({new_n1256_, new_n6235_})
2'b01 : new_n6292_ = 1'b1;
default : new_n6292_ = 1'b0;
endcase
casez ({new_n6285_, new_n6288_})
2'b11 : new_n6293_ = 1'b1;
default : new_n6293_ = 1'b0;
endcase
casez ({new_n2911_, new_n6292_})
2'b01 : new_n6294_ = 1'b1;
default : new_n6294_ = 1'b0;
endcase
casez ({new_n2493_, new_n6293_})
2'b01 : new_n6295_ = 1'b1;
default : new_n6295_ = 1'b0;
endcase
end
endmodule
